`timescale 1ns/100ps
//correct read result:
// 000001a9 000003c0 00000237 0000018b 0000034f 000001bf 00000262 0000036a 00000157 0000005f 000002de 00000325 000000ac 00000308 000002bf 00000332 000001d2 000002b1 00000231 000000ca 00000041 0000011c 000003e7 0000033e 00000388 00000042 000000c4 000001a3 00000189 000001b9 00000028 000000eb 000000af 00000286 000000ca 00000142 00000220 000002b9 00000014 000002c1 0000013c 00000321 00000130 00000144 00000305 0000025e 000002f6 000001d7 000001b4 0000015e 0000001c 000000b8 000001f5 000003f7 000002fc 000003f1 00000361 000003d4 0000009b 00000293 00000261 0000036f 000002c2 00000171 00000176 000001a2 0000003e 00000209 00000259 00000384 000003e0 00000338 00000314 000001b8 00000325 00000163 0000000e 000001ed 000000db 00000224 000000bd 00000327 00000367 00000130 000003ed 00000233 0000036c 000003f8 0000033a 000001eb 00000052 000000ea 0000027f 000002b0 0000012f 00000107 000003c2 0000003c 00000053 0000034b 00000059 00000318 000001f8 000003d5 000000b5 0000026a 000002f5 0000000a 000003fd 00000350 00000304 00000070 00000379 000003d4 00000366 00000189 00000040 00000028 00000130 000002e0 00000105 000000d0 00000058 0000034e 00000154 00000279 0000018b 00000182 00000317 00000365 000000f1 0000010b 000000a5 00000331 00000266 000003f9 000000ca 000000bb 0000017d 00000141 00000371 000000d9 000003f0 00000328 000001e6 00000159 000000a4 000001c5 00000125 000001a1 000001a1 00000311 000000dd 000002f7 0000001f 0000038b 0000028b 000002dc 00000094 00000101 00000074 000000dd 000003ef 000003af 000003fc 00000354 000000e4 00000140 0000008e 00000106 00000011 000001f1 0000036a 00000004 000002e0 0000003a 00000224 000001dc 00000018 00000088 000003ce 0000005a 000003ef 00000171 00000134 000002ac 000003dc 000000b1 000002e6 0000006e 0000034d 000001cb 000000e2 0000003e 0000035d 0000008e 00000289 000003bb 000003a3 00000391 00000395 000003be 0000028d 0000022c 000003ca 000002e2 0000000e 000002ac 0000031f 00000105 000001c1 00000361 000002bd 00000314 0000026d 0000025d 000003ea 0000005c 000001f1 000002fb 000002d1 000001c0 00000344 000002fa 0000022e 000000d3 00000271 00000383 00000050 000002d6 0000014f 000003be 00000198 000000fe 0000036a 00000088 000001b2 00000147 000001a7 000001ca 00000045 00000391 0000030d 000001b3 0000018c 0000033e 00000114 0000036e 000001e3 00000177 000000a0 00000153 0000039f 000000ce 00000291 000002c5

module cache_tb();

`define DATA_COUNT (256)
`define RDWR_COUNT (6*`DATA_COUNT)

reg wr_cycle           [`RDWR_COUNT];
reg rd_cycle           [`RDWR_COUNT];
reg [31:0] addr_rom    [`RDWR_COUNT];
reg [31:0] wr_data_rom [`RDWR_COUNT];
reg [31:0] validation_data [`DATA_COUNT];

initial begin
    // 256 sequence write cycles
    rd_cycle[    0] = 1'b0;  wr_cycle[    0] = 1'b1;  addr_rom[    0]='h00000000;  wr_data_rom[    0]='h00000151;
    rd_cycle[    1] = 1'b0;  wr_cycle[    1] = 1'b1;  addr_rom[    1]='h00000004;  wr_data_rom[    1]='h0000030a;
    rd_cycle[    2] = 1'b0;  wr_cycle[    2] = 1'b1;  addr_rom[    2]='h00000008;  wr_data_rom[    2]='h00000101;
    rd_cycle[    3] = 1'b0;  wr_cycle[    3] = 1'b1;  addr_rom[    3]='h0000000c;  wr_data_rom[    3]='h00000183;
    rd_cycle[    4] = 1'b0;  wr_cycle[    4] = 1'b1;  addr_rom[    4]='h00000010;  wr_data_rom[    4]='h000001b3;
    rd_cycle[    5] = 1'b0;  wr_cycle[    5] = 1'b1;  addr_rom[    5]='h00000014;  wr_data_rom[    5]='h00000161;
    rd_cycle[    6] = 1'b0;  wr_cycle[    6] = 1'b1;  addr_rom[    6]='h00000018;  wr_data_rom[    6]='h0000004f;
    rd_cycle[    7] = 1'b0;  wr_cycle[    7] = 1'b1;  addr_rom[    7]='h0000001c;  wr_data_rom[    7]='h0000036a;
    rd_cycle[    8] = 1'b0;  wr_cycle[    8] = 1'b1;  addr_rom[    8]='h00000020;  wr_data_rom[    8]='h0000016c;
    rd_cycle[    9] = 1'b0;  wr_cycle[    9] = 1'b1;  addr_rom[    9]='h00000024;  wr_data_rom[    9]='h00000217;
    rd_cycle[   10] = 1'b0;  wr_cycle[   10] = 1'b1;  addr_rom[   10]='h00000028;  wr_data_rom[   10]='h000002de;
    rd_cycle[   11] = 1'b0;  wr_cycle[   11] = 1'b1;  addr_rom[   11]='h0000002c;  wr_data_rom[   11]='h00000325;
    rd_cycle[   12] = 1'b0;  wr_cycle[   12] = 1'b1;  addr_rom[   12]='h00000030;  wr_data_rom[   12]='h000001e3;
    rd_cycle[   13] = 1'b0;  wr_cycle[   13] = 1'b1;  addr_rom[   13]='h00000034;  wr_data_rom[   13]='h00000388;
    rd_cycle[   14] = 1'b0;  wr_cycle[   14] = 1'b1;  addr_rom[   14]='h00000038;  wr_data_rom[   14]='h000002bf;
    rd_cycle[   15] = 1'b0;  wr_cycle[   15] = 1'b1;  addr_rom[   15]='h0000003c;  wr_data_rom[   15]='h00000197;
    rd_cycle[   16] = 1'b0;  wr_cycle[   16] = 1'b1;  addr_rom[   16]='h00000040;  wr_data_rom[   16]='h000001fd;
    rd_cycle[   17] = 1'b0;  wr_cycle[   17] = 1'b1;  addr_rom[   17]='h00000044;  wr_data_rom[   17]='h000002b1;
    rd_cycle[   18] = 1'b0;  wr_cycle[   18] = 1'b1;  addr_rom[   18]='h00000048;  wr_data_rom[   18]='h000002bf;
    rd_cycle[   19] = 1'b0;  wr_cycle[   19] = 1'b1;  addr_rom[   19]='h0000004c;  wr_data_rom[   19]='h000000ca;
    rd_cycle[   20] = 1'b0;  wr_cycle[   20] = 1'b1;  addr_rom[   20]='h00000050;  wr_data_rom[   20]='h00000341;
    rd_cycle[   21] = 1'b0;  wr_cycle[   21] = 1'b1;  addr_rom[   21]='h00000054;  wr_data_rom[   21]='h0000011c;
    rd_cycle[   22] = 1'b0;  wr_cycle[   22] = 1'b1;  addr_rom[   22]='h00000058;  wr_data_rom[   22]='h000003e7;
    rd_cycle[   23] = 1'b0;  wr_cycle[   23] = 1'b1;  addr_rom[   23]='h0000005c;  wr_data_rom[   23]='h000002f7;
    rd_cycle[   24] = 1'b0;  wr_cycle[   24] = 1'b1;  addr_rom[   24]='h00000060;  wr_data_rom[   24]='h00000225;
    rd_cycle[   25] = 1'b0;  wr_cycle[   25] = 1'b1;  addr_rom[   25]='h00000064;  wr_data_rom[   25]='h0000015f;
    rd_cycle[   26] = 1'b0;  wr_cycle[   26] = 1'b1;  addr_rom[   26]='h00000068;  wr_data_rom[   26]='h000000c4;
    rd_cycle[   27] = 1'b0;  wr_cycle[   27] = 1'b1;  addr_rom[   27]='h0000006c;  wr_data_rom[   27]='h000001a3;
    rd_cycle[   28] = 1'b0;  wr_cycle[   28] = 1'b1;  addr_rom[   28]='h00000070;  wr_data_rom[   28]='h00000189;
    rd_cycle[   29] = 1'b0;  wr_cycle[   29] = 1'b1;  addr_rom[   29]='h00000074;  wr_data_rom[   29]='h000003ed;
    rd_cycle[   30] = 1'b0;  wr_cycle[   30] = 1'b1;  addr_rom[   30]='h00000078;  wr_data_rom[   30]='h00000287;
    rd_cycle[   31] = 1'b0;  wr_cycle[   31] = 1'b1;  addr_rom[   31]='h0000007c;  wr_data_rom[   31]='h0000022a;
    rd_cycle[   32] = 1'b0;  wr_cycle[   32] = 1'b1;  addr_rom[   32]='h00000080;  wr_data_rom[   32]='h00000276;
    rd_cycle[   33] = 1'b0;  wr_cycle[   33] = 1'b1;  addr_rom[   33]='h00000084;  wr_data_rom[   33]='h00000175;
    rd_cycle[   34] = 1'b0;  wr_cycle[   34] = 1'b1;  addr_rom[   34]='h00000088;  wr_data_rom[   34]='h0000023b;
    rd_cycle[   35] = 1'b0;  wr_cycle[   35] = 1'b1;  addr_rom[   35]='h0000008c;  wr_data_rom[   35]='h0000015b;
    rd_cycle[   36] = 1'b0;  wr_cycle[   36] = 1'b1;  addr_rom[   36]='h00000090;  wr_data_rom[   36]='h000001a9;
    rd_cycle[   37] = 1'b0;  wr_cycle[   37] = 1'b1;  addr_rom[   37]='h00000094;  wr_data_rom[   37]='h00000125;
    rd_cycle[   38] = 1'b0;  wr_cycle[   38] = 1'b1;  addr_rom[   38]='h00000098;  wr_data_rom[   38]='h000002cd;
    rd_cycle[   39] = 1'b0;  wr_cycle[   39] = 1'b1;  addr_rom[   39]='h0000009c;  wr_data_rom[   39]='h000003ad;
    rd_cycle[   40] = 1'b0;  wr_cycle[   40] = 1'b1;  addr_rom[   40]='h000000a0;  wr_data_rom[   40]='h000003a0;
    rd_cycle[   41] = 1'b0;  wr_cycle[   41] = 1'b1;  addr_rom[   41]='h000000a4;  wr_data_rom[   41]='h00000131;
    rd_cycle[   42] = 1'b0;  wr_cycle[   42] = 1'b1;  addr_rom[   42]='h000000a8;  wr_data_rom[   42]='h00000077;
    rd_cycle[   43] = 1'b0;  wr_cycle[   43] = 1'b1;  addr_rom[   43]='h000000ac;  wr_data_rom[   43]='h00000144;
    rd_cycle[   44] = 1'b0;  wr_cycle[   44] = 1'b1;  addr_rom[   44]='h000000b0;  wr_data_rom[   44]='h000003c5;
    rd_cycle[   45] = 1'b0;  wr_cycle[   45] = 1'b1;  addr_rom[   45]='h000000b4;  wr_data_rom[   45]='h000002e9;
    rd_cycle[   46] = 1'b0;  wr_cycle[   46] = 1'b1;  addr_rom[   46]='h000000b8;  wr_data_rom[   46]='h000001ab;
    rd_cycle[   47] = 1'b0;  wr_cycle[   47] = 1'b1;  addr_rom[   47]='h000000bc;  wr_data_rom[   47]='h00000320;
    rd_cycle[   48] = 1'b0;  wr_cycle[   48] = 1'b1;  addr_rom[   48]='h000000c0;  wr_data_rom[   48]='h000001b4;
    rd_cycle[   49] = 1'b0;  wr_cycle[   49] = 1'b1;  addr_rom[   49]='h000000c4;  wr_data_rom[   49]='h0000015e;
    rd_cycle[   50] = 1'b0;  wr_cycle[   50] = 1'b1;  addr_rom[   50]='h000000c8;  wr_data_rom[   50]='h00000072;
    rd_cycle[   51] = 1'b0;  wr_cycle[   51] = 1'b1;  addr_rom[   51]='h000000cc;  wr_data_rom[   51]='h00000236;
    rd_cycle[   52] = 1'b0;  wr_cycle[   52] = 1'b1;  addr_rom[   52]='h000000d0;  wr_data_rom[   52]='h00000393;
    rd_cycle[   53] = 1'b0;  wr_cycle[   53] = 1'b1;  addr_rom[   53]='h000000d4;  wr_data_rom[   53]='h000003f7;
    rd_cycle[   54] = 1'b0;  wr_cycle[   54] = 1'b1;  addr_rom[   54]='h000000d8;  wr_data_rom[   54]='h000002fc;
    rd_cycle[   55] = 1'b0;  wr_cycle[   55] = 1'b1;  addr_rom[   55]='h000000dc;  wr_data_rom[   55]='h000000eb;
    rd_cycle[   56] = 1'b0;  wr_cycle[   56] = 1'b1;  addr_rom[   56]='h000000e0;  wr_data_rom[   56]='h00000128;
    rd_cycle[   57] = 1'b0;  wr_cycle[   57] = 1'b1;  addr_rom[   57]='h000000e4;  wr_data_rom[   57]='h00000180;
    rd_cycle[   58] = 1'b0;  wr_cycle[   58] = 1'b1;  addr_rom[   58]='h000000e8;  wr_data_rom[   58]='h000000d6;
    rd_cycle[   59] = 1'b0;  wr_cycle[   59] = 1'b1;  addr_rom[   59]='h000000ec;  wr_data_rom[   59]='h000000b4;
    rd_cycle[   60] = 1'b0;  wr_cycle[   60] = 1'b1;  addr_rom[   60]='h000000f0;  wr_data_rom[   60]='h000000f0;
    rd_cycle[   61] = 1'b0;  wr_cycle[   61] = 1'b1;  addr_rom[   61]='h000000f4;  wr_data_rom[   61]='h000003c7;
    rd_cycle[   62] = 1'b0;  wr_cycle[   62] = 1'b1;  addr_rom[   62]='h000000f8;  wr_data_rom[   62]='h00000075;
    rd_cycle[   63] = 1'b0;  wr_cycle[   63] = 1'b1;  addr_rom[   63]='h000000fc;  wr_data_rom[   63]='h000002ee;
    rd_cycle[   64] = 1'b0;  wr_cycle[   64] = 1'b1;  addr_rom[   64]='h00000100;  wr_data_rom[   64]='h000001e1;
    rd_cycle[   65] = 1'b0;  wr_cycle[   65] = 1'b1;  addr_rom[   65]='h00000104;  wr_data_rom[   65]='h000000e1;
    rd_cycle[   66] = 1'b0;  wr_cycle[   66] = 1'b1;  addr_rom[   66]='h00000108;  wr_data_rom[   66]='h000001a1;
    rd_cycle[   67] = 1'b0;  wr_cycle[   67] = 1'b1;  addr_rom[   67]='h0000010c;  wr_data_rom[   67]='h000003a2;
    rd_cycle[   68] = 1'b0;  wr_cycle[   68] = 1'b1;  addr_rom[   68]='h00000110;  wr_data_rom[   68]='h00000065;
    rd_cycle[   69] = 1'b0;  wr_cycle[   69] = 1'b1;  addr_rom[   69]='h00000114;  wr_data_rom[   69]='h00000133;
    rd_cycle[   70] = 1'b0;  wr_cycle[   70] = 1'b1;  addr_rom[   70]='h00000118;  wr_data_rom[   70]='h0000031f;
    rd_cycle[   71] = 1'b0;  wr_cycle[   71] = 1'b1;  addr_rom[   71]='h0000011c;  wr_data_rom[   71]='h00000338;
    rd_cycle[   72] = 1'b0;  wr_cycle[   72] = 1'b1;  addr_rom[   72]='h00000120;  wr_data_rom[   72]='h0000034d;
    rd_cycle[   73] = 1'b0;  wr_cycle[   73] = 1'b1;  addr_rom[   73]='h00000124;  wr_data_rom[   73]='h000003c2;
    rd_cycle[   74] = 1'b0;  wr_cycle[   74] = 1'b1;  addr_rom[   74]='h00000128;  wr_data_rom[   74]='h0000007f;
    rd_cycle[   75] = 1'b0;  wr_cycle[   75] = 1'b1;  addr_rom[   75]='h0000012c;  wr_data_rom[   75]='h0000008f;
    rd_cycle[   76] = 1'b0;  wr_cycle[   76] = 1'b1;  addr_rom[   76]='h00000130;  wr_data_rom[   76]='h00000267;
    rd_cycle[   77] = 1'b0;  wr_cycle[   77] = 1'b1;  addr_rom[   77]='h00000134;  wr_data_rom[   77]='h000001ed;
    rd_cycle[   78] = 1'b0;  wr_cycle[   78] = 1'b1;  addr_rom[   78]='h00000138;  wr_data_rom[   78]='h0000007d;
    rd_cycle[   79] = 1'b0;  wr_cycle[   79] = 1'b1;  addr_rom[   79]='h0000013c;  wr_data_rom[   79]='h000001a0;
    rd_cycle[   80] = 1'b0;  wr_cycle[   80] = 1'b1;  addr_rom[   80]='h00000140;  wr_data_rom[   80]='h000000e8;
    rd_cycle[   81] = 1'b0;  wr_cycle[   81] = 1'b1;  addr_rom[   81]='h00000144;  wr_data_rom[   81]='h00000031;
    rd_cycle[   82] = 1'b0;  wr_cycle[   82] = 1'b1;  addr_rom[   82]='h00000148;  wr_data_rom[   82]='h00000237;
    rd_cycle[   83] = 1'b0;  wr_cycle[   83] = 1'b1;  addr_rom[   83]='h0000014c;  wr_data_rom[   83]='h0000034b;
    rd_cycle[   84] = 1'b0;  wr_cycle[   84] = 1'b1;  addr_rom[   84]='h00000150;  wr_data_rom[   84]='h000003ed;
    rd_cycle[   85] = 1'b0;  wr_cycle[   85] = 1'b1;  addr_rom[   85]='h00000154;  wr_data_rom[   85]='h00000363;
    rd_cycle[   86] = 1'b0;  wr_cycle[   86] = 1'b1;  addr_rom[   86]='h00000158;  wr_data_rom[   86]='h000003d1;
    rd_cycle[   87] = 1'b0;  wr_cycle[   87] = 1'b1;  addr_rom[   87]='h0000015c;  wr_data_rom[   87]='h00000250;
    rd_cycle[   88] = 1'b0;  wr_cycle[   88] = 1'b1;  addr_rom[   88]='h00000160;  wr_data_rom[   88]='h00000396;
    rd_cycle[   89] = 1'b0;  wr_cycle[   89] = 1'b1;  addr_rom[   89]='h00000164;  wr_data_rom[   89]='h0000014c;
    rd_cycle[   90] = 1'b0;  wr_cycle[   90] = 1'b1;  addr_rom[   90]='h00000168;  wr_data_rom[   90]='h00000030;
    rd_cycle[   91] = 1'b0;  wr_cycle[   91] = 1'b1;  addr_rom[   91]='h0000016c;  wr_data_rom[   91]='h000002fe;
    rd_cycle[   92] = 1'b0;  wr_cycle[   92] = 1'b1;  addr_rom[   92]='h00000170;  wr_data_rom[   92]='h0000027f;
    rd_cycle[   93] = 1'b0;  wr_cycle[   93] = 1'b1;  addr_rom[   93]='h00000174;  wr_data_rom[   93]='h000003bf;
    rd_cycle[   94] = 1'b0;  wr_cycle[   94] = 1'b1;  addr_rom[   94]='h00000178;  wr_data_rom[   94]='h0000038b;
    rd_cycle[   95] = 1'b0;  wr_cycle[   95] = 1'b1;  addr_rom[   95]='h0000017c;  wr_data_rom[   95]='h00000107;
    rd_cycle[   96] = 1'b0;  wr_cycle[   96] = 1'b1;  addr_rom[   96]='h00000180;  wr_data_rom[   96]='h00000016;
    rd_cycle[   97] = 1'b0;  wr_cycle[   97] = 1'b1;  addr_rom[   97]='h00000184;  wr_data_rom[   97]='h0000003c;
    rd_cycle[   98] = 1'b0;  wr_cycle[   98] = 1'b1;  addr_rom[   98]='h00000188;  wr_data_rom[   98]='h0000003d;
    rd_cycle[   99] = 1'b0;  wr_cycle[   99] = 1'b1;  addr_rom[   99]='h0000018c;  wr_data_rom[   99]='h00000230;
    rd_cycle[  100] = 1'b0;  wr_cycle[  100] = 1'b1;  addr_rom[  100]='h00000190;  wr_data_rom[  100]='h00000276;
    rd_cycle[  101] = 1'b0;  wr_cycle[  101] = 1'b1;  addr_rom[  101]='h00000194;  wr_data_rom[  101]='h00000318;
    rd_cycle[  102] = 1'b0;  wr_cycle[  102] = 1'b1;  addr_rom[  102]='h00000198;  wr_data_rom[  102]='h000002de;
    rd_cycle[  103] = 1'b0;  wr_cycle[  103] = 1'b1;  addr_rom[  103]='h0000019c;  wr_data_rom[  103]='h000003cc;
    rd_cycle[  104] = 1'b0;  wr_cycle[  104] = 1'b1;  addr_rom[  104]='h000001a0;  wr_data_rom[  104]='h00000266;
    rd_cycle[  105] = 1'b0;  wr_cycle[  105] = 1'b1;  addr_rom[  105]='h000001a4;  wr_data_rom[  105]='h00000150;
    rd_cycle[  106] = 1'b0;  wr_cycle[  106] = 1'b1;  addr_rom[  106]='h000001a8;  wr_data_rom[  106]='h000002f5;
    rd_cycle[  107] = 1'b0;  wr_cycle[  107] = 1'b1;  addr_rom[  107]='h000001ac;  wr_data_rom[  107]='h0000000a;
    rd_cycle[  108] = 1'b0;  wr_cycle[  108] = 1'b1;  addr_rom[  108]='h000001b0;  wr_data_rom[  108]='h000001aa;
    rd_cycle[  109] = 1'b0;  wr_cycle[  109] = 1'b1;  addr_rom[  109]='h000001b4;  wr_data_rom[  109]='h00000350;
    rd_cycle[  110] = 1'b0;  wr_cycle[  110] = 1'b1;  addr_rom[  110]='h000001b8;  wr_data_rom[  110]='h000000ac;
    rd_cycle[  111] = 1'b0;  wr_cycle[  111] = 1'b1;  addr_rom[  111]='h000001bc;  wr_data_rom[  111]='h0000029a;
    rd_cycle[  112] = 1'b0;  wr_cycle[  112] = 1'b1;  addr_rom[  112]='h000001c0;  wr_data_rom[  112]='h00000052;
    rd_cycle[  113] = 1'b0;  wr_cycle[  113] = 1'b1;  addr_rom[  113]='h000001c4;  wr_data_rom[  113]='h000003d4;
    rd_cycle[  114] = 1'b0;  wr_cycle[  114] = 1'b1;  addr_rom[  114]='h000001c8;  wr_data_rom[  114]='h000001dd;
    rd_cycle[  115] = 1'b0;  wr_cycle[  115] = 1'b1;  addr_rom[  115]='h000001cc;  wr_data_rom[  115]='h00000179;
    rd_cycle[  116] = 1'b0;  wr_cycle[  116] = 1'b1;  addr_rom[  116]='h000001d0;  wr_data_rom[  116]='h00000216;
    rd_cycle[  117] = 1'b0;  wr_cycle[  117] = 1'b1;  addr_rom[  117]='h000001d4;  wr_data_rom[  117]='h00000394;
    rd_cycle[  118] = 1'b0;  wr_cycle[  118] = 1'b1;  addr_rom[  118]='h000001d8;  wr_data_rom[  118]='h00000130;
    rd_cycle[  119] = 1'b0;  wr_cycle[  119] = 1'b1;  addr_rom[  119]='h000001dc;  wr_data_rom[  119]='h000000c3;
    rd_cycle[  120] = 1'b0;  wr_cycle[  120] = 1'b1;  addr_rom[  120]='h000001e0;  wr_data_rom[  120]='h0000017b;
    rd_cycle[  121] = 1'b0;  wr_cycle[  121] = 1'b1;  addr_rom[  121]='h000001e4;  wr_data_rom[  121]='h000002fa;
    rd_cycle[  122] = 1'b0;  wr_cycle[  122] = 1'b1;  addr_rom[  122]='h000001e8;  wr_data_rom[  122]='h0000014e;
    rd_cycle[  123] = 1'b0;  wr_cycle[  123] = 1'b1;  addr_rom[  123]='h000001ec;  wr_data_rom[  123]='h000000eb;
    rd_cycle[  124] = 1'b0;  wr_cycle[  124] = 1'b1;  addr_rom[  124]='h000001f0;  wr_data_rom[  124]='h00000154;
    rd_cycle[  125] = 1'b0;  wr_cycle[  125] = 1'b1;  addr_rom[  125]='h000001f4;  wr_data_rom[  125]='h000001fc;
    rd_cycle[  126] = 1'b0;  wr_cycle[  126] = 1'b1;  addr_rom[  126]='h000001f8;  wr_data_rom[  126]='h000001d9;
    rd_cycle[  127] = 1'b0;  wr_cycle[  127] = 1'b1;  addr_rom[  127]='h000001fc;  wr_data_rom[  127]='h000003ac;
    rd_cycle[  128] = 1'b0;  wr_cycle[  128] = 1'b1;  addr_rom[  128]='h00000200;  wr_data_rom[  128]='h00000317;
    rd_cycle[  129] = 1'b0;  wr_cycle[  129] = 1'b1;  addr_rom[  129]='h00000204;  wr_data_rom[  129]='h00000365;
    rd_cycle[  130] = 1'b0;  wr_cycle[  130] = 1'b1;  addr_rom[  130]='h00000208;  wr_data_rom[  130]='h000000f1;
    rd_cycle[  131] = 1'b0;  wr_cycle[  131] = 1'b1;  addr_rom[  131]='h0000020c;  wr_data_rom[  131]='h000003ec;
    rd_cycle[  132] = 1'b0;  wr_cycle[  132] = 1'b1;  addr_rom[  132]='h00000210;  wr_data_rom[  132]='h0000005c;
    rd_cycle[  133] = 1'b0;  wr_cycle[  133] = 1'b1;  addr_rom[  133]='h00000214;  wr_data_rom[  133]='h00000331;
    rd_cycle[  134] = 1'b0;  wr_cycle[  134] = 1'b1;  addr_rom[  134]='h00000218;  wr_data_rom[  134]='h00000359;
    rd_cycle[  135] = 1'b0;  wr_cycle[  135] = 1'b1;  addr_rom[  135]='h0000021c;  wr_data_rom[  135]='h000001d4;
    rd_cycle[  136] = 1'b0;  wr_cycle[  136] = 1'b1;  addr_rom[  136]='h00000220;  wr_data_rom[  136]='h00000308;
    rd_cycle[  137] = 1'b0;  wr_cycle[  137] = 1'b1;  addr_rom[  137]='h00000224;  wr_data_rom[  137]='h000000bb;
    rd_cycle[  138] = 1'b0;  wr_cycle[  138] = 1'b1;  addr_rom[  138]='h00000228;  wr_data_rom[  138]='h00000151;
    rd_cycle[  139] = 1'b0;  wr_cycle[  139] = 1'b1;  addr_rom[  139]='h0000022c;  wr_data_rom[  139]='h000003c5;
    rd_cycle[  140] = 1'b0;  wr_cycle[  140] = 1'b1;  addr_rom[  140]='h00000230;  wr_data_rom[  140]='h00000371;
    rd_cycle[  141] = 1'b0;  wr_cycle[  141] = 1'b1;  addr_rom[  141]='h00000234;  wr_data_rom[  141]='h000002ce;
    rd_cycle[  142] = 1'b0;  wr_cycle[  142] = 1'b1;  addr_rom[  142]='h00000238;  wr_data_rom[  142]='h000001ef;
    rd_cycle[  143] = 1'b0;  wr_cycle[  143] = 1'b1;  addr_rom[  143]='h0000023c;  wr_data_rom[  143]='h00000328;
    rd_cycle[  144] = 1'b0;  wr_cycle[  144] = 1'b1;  addr_rom[  144]='h00000240;  wr_data_rom[  144]='h000001e6;
    rd_cycle[  145] = 1'b0;  wr_cycle[  145] = 1'b1;  addr_rom[  145]='h00000244;  wr_data_rom[  145]='h00000169;
    rd_cycle[  146] = 1'b0;  wr_cycle[  146] = 1'b1;  addr_rom[  146]='h00000248;  wr_data_rom[  146]='h0000023e;
    rd_cycle[  147] = 1'b0;  wr_cycle[  147] = 1'b1;  addr_rom[  147]='h0000024c;  wr_data_rom[  147]='h00000368;
    rd_cycle[  148] = 1'b0;  wr_cycle[  148] = 1'b1;  addr_rom[  148]='h00000250;  wr_data_rom[  148]='h000003e0;
    rd_cycle[  149] = 1'b0;  wr_cycle[  149] = 1'b1;  addr_rom[  149]='h00000254;  wr_data_rom[  149]='h00000084;
    rd_cycle[  150] = 1'b0;  wr_cycle[  150] = 1'b1;  addr_rom[  150]='h00000258;  wr_data_rom[  150]='h0000027f;
    rd_cycle[  151] = 1'b0;  wr_cycle[  151] = 1'b1;  addr_rom[  151]='h0000025c;  wr_data_rom[  151]='h00000311;
    rd_cycle[  152] = 1'b0;  wr_cycle[  152] = 1'b1;  addr_rom[  152]='h00000260;  wr_data_rom[  152]='h000002b9;
    rd_cycle[  153] = 1'b0;  wr_cycle[  153] = 1'b1;  addr_rom[  153]='h00000264;  wr_data_rom[  153]='h00000134;
    rd_cycle[  154] = 1'b0;  wr_cycle[  154] = 1'b1;  addr_rom[  154]='h00000268;  wr_data_rom[  154]='h00000138;
    rd_cycle[  155] = 1'b0;  wr_cycle[  155] = 1'b1;  addr_rom[  155]='h0000026c;  wr_data_rom[  155]='h00000071;
    rd_cycle[  156] = 1'b0;  wr_cycle[  156] = 1'b1;  addr_rom[  156]='h00000270;  wr_data_rom[  156]='h0000028b;
    rd_cycle[  157] = 1'b0;  wr_cycle[  157] = 1'b1;  addr_rom[  157]='h00000274;  wr_data_rom[  157]='h00000278;
    rd_cycle[  158] = 1'b0;  wr_cycle[  158] = 1'b1;  addr_rom[  158]='h00000278;  wr_data_rom[  158]='h00000234;
    rd_cycle[  159] = 1'b0;  wr_cycle[  159] = 1'b1;  addr_rom[  159]='h0000027c;  wr_data_rom[  159]='h00000101;
    rd_cycle[  160] = 1'b0;  wr_cycle[  160] = 1'b1;  addr_rom[  160]='h00000280;  wr_data_rom[  160]='h0000027c;
    rd_cycle[  161] = 1'b0;  wr_cycle[  161] = 1'b1;  addr_rom[  161]='h00000284;  wr_data_rom[  161]='h000000dd;
    rd_cycle[  162] = 1'b0;  wr_cycle[  162] = 1'b1;  addr_rom[  162]='h00000288;  wr_data_rom[  162]='h0000031d;
    rd_cycle[  163] = 1'b0;  wr_cycle[  163] = 1'b1;  addr_rom[  163]='h0000028c;  wr_data_rom[  163]='h000002a6;
    rd_cycle[  164] = 1'b0;  wr_cycle[  164] = 1'b1;  addr_rom[  164]='h00000290;  wr_data_rom[  164]='h000003fc;
    rd_cycle[  165] = 1'b0;  wr_cycle[  165] = 1'b1;  addr_rom[  165]='h00000294;  wr_data_rom[  165]='h00000142;
    rd_cycle[  166] = 1'b0;  wr_cycle[  166] = 1'b1;  addr_rom[  166]='h00000298;  wr_data_rom[  166]='h000001e6;
    rd_cycle[  167] = 1'b0;  wr_cycle[  167] = 1'b1;  addr_rom[  167]='h0000029c;  wr_data_rom[  167]='h00000387;
    rd_cycle[  168] = 1'b0;  wr_cycle[  168] = 1'b1;  addr_rom[  168]='h000002a0;  wr_data_rom[  168]='h00000140;
    rd_cycle[  169] = 1'b0;  wr_cycle[  169] = 1'b1;  addr_rom[  169]='h000002a4;  wr_data_rom[  169]='h000002b6;
    rd_cycle[  170] = 1'b0;  wr_cycle[  170] = 1'b1;  addr_rom[  170]='h000002a8;  wr_data_rom[  170]='h0000027f;
    rd_cycle[  171] = 1'b0;  wr_cycle[  171] = 1'b1;  addr_rom[  171]='h000002ac;  wr_data_rom[  171]='h00000131;
    rd_cycle[  172] = 1'b0;  wr_cycle[  172] = 1'b1;  addr_rom[  172]='h000002b0;  wr_data_rom[  172]='h0000036a;
    rd_cycle[  173] = 1'b0;  wr_cycle[  173] = 1'b1;  addr_rom[  173]='h000002b4;  wr_data_rom[  173]='h00000190;
    rd_cycle[  174] = 1'b0;  wr_cycle[  174] = 1'b1;  addr_rom[  174]='h000002b8;  wr_data_rom[  174]='h000001d5;
    rd_cycle[  175] = 1'b0;  wr_cycle[  175] = 1'b1;  addr_rom[  175]='h000002bc;  wr_data_rom[  175]='h0000003a;
    rd_cycle[  176] = 1'b0;  wr_cycle[  176] = 1'b1;  addr_rom[  176]='h000002c0;  wr_data_rom[  176]='h000000b6;
    rd_cycle[  177] = 1'b0;  wr_cycle[  177] = 1'b1;  addr_rom[  177]='h000002c4;  wr_data_rom[  177]='h000003f1;
    rd_cycle[  178] = 1'b0;  wr_cycle[  178] = 1'b1;  addr_rom[  178]='h000002c8;  wr_data_rom[  178]='h00000082;
    rd_cycle[  179] = 1'b0;  wr_cycle[  179] = 1'b1;  addr_rom[  179]='h000002cc;  wr_data_rom[  179]='h00000268;
    rd_cycle[  180] = 1'b0;  wr_cycle[  180] = 1'b1;  addr_rom[  180]='h000002d0;  wr_data_rom[  180]='h000002b3;
    rd_cycle[  181] = 1'b0;  wr_cycle[  181] = 1'b1;  addr_rom[  181]='h000002d4;  wr_data_rom[  181]='h000003e7;
    rd_cycle[  182] = 1'b0;  wr_cycle[  182] = 1'b1;  addr_rom[  182]='h000002d8;  wr_data_rom[  182]='h0000027e;
    rd_cycle[  183] = 1'b0;  wr_cycle[  183] = 1'b1;  addr_rom[  183]='h000002dc;  wr_data_rom[  183]='h00000171;
    rd_cycle[  184] = 1'b0;  wr_cycle[  184] = 1'b1;  addr_rom[  184]='h000002e0;  wr_data_rom[  184]='h0000003d;
    rd_cycle[  185] = 1'b0;  wr_cycle[  185] = 1'b1;  addr_rom[  185]='h000002e4;  wr_data_rom[  185]='h000003a1;
    rd_cycle[  186] = 1'b0;  wr_cycle[  186] = 1'b1;  addr_rom[  186]='h000002e8;  wr_data_rom[  186]='h000003dc;
    rd_cycle[  187] = 1'b0;  wr_cycle[  187] = 1'b1;  addr_rom[  187]='h000002ec;  wr_data_rom[  187]='h000000b1;
    rd_cycle[  188] = 1'b0;  wr_cycle[  188] = 1'b1;  addr_rom[  188]='h000002f0;  wr_data_rom[  188]='h000002e6;
    rd_cycle[  189] = 1'b0;  wr_cycle[  189] = 1'b1;  addr_rom[  189]='h000002f4;  wr_data_rom[  189]='h0000027a;
    rd_cycle[  190] = 1'b0;  wr_cycle[  190] = 1'b1;  addr_rom[  190]='h000002f8;  wr_data_rom[  190]='h0000034d;
    rd_cycle[  191] = 1'b0;  wr_cycle[  191] = 1'b1;  addr_rom[  191]='h000002fc;  wr_data_rom[  191]='h000001cb;
    rd_cycle[  192] = 1'b0;  wr_cycle[  192] = 1'b1;  addr_rom[  192]='h00000300;  wr_data_rom[  192]='h000000a0;
    rd_cycle[  193] = 1'b0;  wr_cycle[  193] = 1'b1;  addr_rom[  193]='h00000304;  wr_data_rom[  193]='h0000003e;
    rd_cycle[  194] = 1'b0;  wr_cycle[  194] = 1'b1;  addr_rom[  194]='h00000308;  wr_data_rom[  194]='h00000267;
    rd_cycle[  195] = 1'b0;  wr_cycle[  195] = 1'b1;  addr_rom[  195]='h0000030c;  wr_data_rom[  195]='h000000f9;
    rd_cycle[  196] = 1'b0;  wr_cycle[  196] = 1'b1;  addr_rom[  196]='h00000310;  wr_data_rom[  196]='h00000289;
    rd_cycle[  197] = 1'b0;  wr_cycle[  197] = 1'b1;  addr_rom[  197]='h00000314;  wr_data_rom[  197]='h00000384;
    rd_cycle[  198] = 1'b0;  wr_cycle[  198] = 1'b1;  addr_rom[  198]='h00000318;  wr_data_rom[  198]='h00000033;
    rd_cycle[  199] = 1'b0;  wr_cycle[  199] = 1'b1;  addr_rom[  199]='h0000031c;  wr_data_rom[  199]='h000001b1;
    rd_cycle[  200] = 1'b0;  wr_cycle[  200] = 1'b1;  addr_rom[  200]='h00000320;  wr_data_rom[  200]='h00000304;
    rd_cycle[  201] = 1'b0;  wr_cycle[  201] = 1'b1;  addr_rom[  201]='h00000324;  wr_data_rom[  201]='h000002eb;
    rd_cycle[  202] = 1'b0;  wr_cycle[  202] = 1'b1;  addr_rom[  202]='h00000328;  wr_data_rom[  202]='h0000028d;
    rd_cycle[  203] = 1'b0;  wr_cycle[  203] = 1'b1;  addr_rom[  203]='h0000032c;  wr_data_rom[  203]='h00000093;
    rd_cycle[  204] = 1'b0;  wr_cycle[  204] = 1'b1;  addr_rom[  204]='h00000330;  wr_data_rom[  204]='h000001c3;
    rd_cycle[  205] = 1'b0;  wr_cycle[  205] = 1'b1;  addr_rom[  205]='h00000334;  wr_data_rom[  205]='h00000226;
    rd_cycle[  206] = 1'b0;  wr_cycle[  206] = 1'b1;  addr_rom[  206]='h00000338;  wr_data_rom[  206]='h0000000e;
    rd_cycle[  207] = 1'b0;  wr_cycle[  207] = 1'b1;  addr_rom[  207]='h0000033c;  wr_data_rom[  207]='h000002ac;
    rd_cycle[  208] = 1'b0;  wr_cycle[  208] = 1'b1;  addr_rom[  208]='h00000340;  wr_data_rom[  208]='h0000011b;
    rd_cycle[  209] = 1'b0;  wr_cycle[  209] = 1'b1;  addr_rom[  209]='h00000344;  wr_data_rom[  209]='h00000359;
    rd_cycle[  210] = 1'b0;  wr_cycle[  210] = 1'b1;  addr_rom[  210]='h00000348;  wr_data_rom[  210]='h00000091;
    rd_cycle[  211] = 1'b0;  wr_cycle[  211] = 1'b1;  addr_rom[  211]='h0000034c;  wr_data_rom[  211]='h00000021;
    rd_cycle[  212] = 1'b0;  wr_cycle[  212] = 1'b1;  addr_rom[  212]='h00000350;  wr_data_rom[  212]='h000002bd;
    rd_cycle[  213] = 1'b0;  wr_cycle[  213] = 1'b1;  addr_rom[  213]='h00000354;  wr_data_rom[  213]='h00000314;
    rd_cycle[  214] = 1'b0;  wr_cycle[  214] = 1'b1;  addr_rom[  214]='h00000358;  wr_data_rom[  214]='h0000032b;
    rd_cycle[  215] = 1'b0;  wr_cycle[  215] = 1'b1;  addr_rom[  215]='h0000035c;  wr_data_rom[  215]='h0000025d;
    rd_cycle[  216] = 1'b0;  wr_cycle[  216] = 1'b1;  addr_rom[  216]='h00000360;  wr_data_rom[  216]='h0000036a;
    rd_cycle[  217] = 1'b0;  wr_cycle[  217] = 1'b1;  addr_rom[  217]='h00000364;  wr_data_rom[  217]='h000001c0;
    rd_cycle[  218] = 1'b0;  wr_cycle[  218] = 1'b1;  addr_rom[  218]='h00000368;  wr_data_rom[  218]='h0000014d;
    rd_cycle[  219] = 1'b0;  wr_cycle[  219] = 1'b1;  addr_rom[  219]='h0000036c;  wr_data_rom[  219]='h0000032f;
    rd_cycle[  220] = 1'b0;  wr_cycle[  220] = 1'b1;  addr_rom[  220]='h00000370;  wr_data_rom[  220]='h00000332;
    rd_cycle[  221] = 1'b0;  wr_cycle[  221] = 1'b1;  addr_rom[  221]='h00000374;  wr_data_rom[  221]='h000001c0;
    rd_cycle[  222] = 1'b0;  wr_cycle[  222] = 1'b1;  addr_rom[  222]='h00000378;  wr_data_rom[  222]='h0000019b;
    rd_cycle[  223] = 1'b0;  wr_cycle[  223] = 1'b1;  addr_rom[  223]='h0000037c;  wr_data_rom[  223]='h00000225;
    rd_cycle[  224] = 1'b0;  wr_cycle[  224] = 1'b1;  addr_rom[  224]='h00000380;  wr_data_rom[  224]='h00000101;
    rd_cycle[  225] = 1'b0;  wr_cycle[  225] = 1'b1;  addr_rom[  225]='h00000384;  wr_data_rom[  225]='h00000080;
    rd_cycle[  226] = 1'b0;  wr_cycle[  226] = 1'b1;  addr_rom[  226]='h00000388;  wr_data_rom[  226]='h00000156;
    rd_cycle[  227] = 1'b0;  wr_cycle[  227] = 1'b1;  addr_rom[  227]='h0000038c;  wr_data_rom[  227]='h000003d6;
    rd_cycle[  228] = 1'b0;  wr_cycle[  228] = 1'b1;  addr_rom[  228]='h00000390;  wr_data_rom[  228]='h000002dc;
    rd_cycle[  229] = 1'b0;  wr_cycle[  229] = 1'b1;  addr_rom[  229]='h00000394;  wr_data_rom[  229]='h000000b5;
    rd_cycle[  230] = 1'b0;  wr_cycle[  230] = 1'b1;  addr_rom[  230]='h00000398;  wr_data_rom[  230]='h000000fa;
    rd_cycle[  231] = 1'b0;  wr_cycle[  231] = 1'b1;  addr_rom[  231]='h0000039c;  wr_data_rom[  231]='h000001f4;
    rd_cycle[  232] = 1'b0;  wr_cycle[  232] = 1'b1;  addr_rom[  232]='h000003a0;  wr_data_rom[  232]='h00000198;
    rd_cycle[  233] = 1'b0;  wr_cycle[  233] = 1'b1;  addr_rom[  233]='h000003a4;  wr_data_rom[  233]='h00000291;
    rd_cycle[  234] = 1'b0;  wr_cycle[  234] = 1'b1;  addr_rom[  234]='h000003a8;  wr_data_rom[  234]='h0000036a;
    rd_cycle[  235] = 1'b0;  wr_cycle[  235] = 1'b1;  addr_rom[  235]='h000003ac;  wr_data_rom[  235]='h00000005;
    rd_cycle[  236] = 1'b0;  wr_cycle[  236] = 1'b1;  addr_rom[  236]='h000003b0;  wr_data_rom[  236]='h000001a1;
    rd_cycle[  237] = 1'b0;  wr_cycle[  237] = 1'b1;  addr_rom[  237]='h000003b4;  wr_data_rom[  237]='h0000035a;
    rd_cycle[  238] = 1'b0;  wr_cycle[  238] = 1'b1;  addr_rom[  238]='h000003b8;  wr_data_rom[  238]='h000000f7;
    rd_cycle[  239] = 1'b0;  wr_cycle[  239] = 1'b1;  addr_rom[  239]='h000003bc;  wr_data_rom[  239]='h000001eb;
    rd_cycle[  240] = 1'b0;  wr_cycle[  240] = 1'b1;  addr_rom[  240]='h000003c0;  wr_data_rom[  240]='h0000021f;
    rd_cycle[  241] = 1'b0;  wr_cycle[  241] = 1'b1;  addr_rom[  241]='h000003c4;  wr_data_rom[  241]='h00000365;
    rd_cycle[  242] = 1'b0;  wr_cycle[  242] = 1'b1;  addr_rom[  242]='h000003c8;  wr_data_rom[  242]='h0000030d;
    rd_cycle[  243] = 1'b0;  wr_cycle[  243] = 1'b1;  addr_rom[  243]='h000003cc;  wr_data_rom[  243]='h000001b3;
    rd_cycle[  244] = 1'b0;  wr_cycle[  244] = 1'b1;  addr_rom[  244]='h000003d0;  wr_data_rom[  244]='h00000278;
    rd_cycle[  245] = 1'b0;  wr_cycle[  245] = 1'b1;  addr_rom[  245]='h000003d4;  wr_data_rom[  245]='h000002ad;
    rd_cycle[  246] = 1'b0;  wr_cycle[  246] = 1'b1;  addr_rom[  246]='h000003d8;  wr_data_rom[  246]='h000002c0;
    rd_cycle[  247] = 1'b0;  wr_cycle[  247] = 1'b1;  addr_rom[  247]='h000003dc;  wr_data_rom[  247]='h0000029d;
    rd_cycle[  248] = 1'b0;  wr_cycle[  248] = 1'b1;  addr_rom[  248]='h000003e0;  wr_data_rom[  248]='h0000024f;
    rd_cycle[  249] = 1'b0;  wr_cycle[  249] = 1'b1;  addr_rom[  249]='h000003e4;  wr_data_rom[  249]='h00000177;
    rd_cycle[  250] = 1'b0;  wr_cycle[  250] = 1'b1;  addr_rom[  250]='h000003e8;  wr_data_rom[  250]='h00000040;
    rd_cycle[  251] = 1'b0;  wr_cycle[  251] = 1'b1;  addr_rom[  251]='h000003ec;  wr_data_rom[  251]='h000003f4;
    rd_cycle[  252] = 1'b0;  wr_cycle[  252] = 1'b1;  addr_rom[  252]='h000003f0;  wr_data_rom[  252]='h0000034c;
    rd_cycle[  253] = 1'b0;  wr_cycle[  253] = 1'b1;  addr_rom[  253]='h000003f4;  wr_data_rom[  253]='h00000400;
    rd_cycle[  254] = 1'b0;  wr_cycle[  254] = 1'b1;  addr_rom[  254]='h000003f8;  wr_data_rom[  254]='h0000039c;
    rd_cycle[  255] = 1'b0;  wr_cycle[  255] = 1'b1;  addr_rom[  255]='h000003fc;  wr_data_rom[  255]='h000002c5;
    // 768 random read and write cycles
    rd_cycle[  256] = 1'b1;  wr_cycle[  256] = 1'b0;  addr_rom[  256]='h00000118;  wr_data_rom[  256]='h00000000;
    rd_cycle[  257] = 1'b0;  wr_cycle[  257] = 1'b1;  addr_rom[  257]='h000001fc;  wr_data_rom[  257]='h000003a3;
    rd_cycle[  258] = 1'b0;  wr_cycle[  258] = 1'b1;  addr_rom[  258]='h00000080;  wr_data_rom[  258]='h00000379;
    rd_cycle[  259] = 1'b1;  wr_cycle[  259] = 1'b0;  addr_rom[  259]='h000002fc;  wr_data_rom[  259]='h00000000;
    rd_cycle[  260] = 1'b0;  wr_cycle[  260] = 1'b1;  addr_rom[  260]='h000003ec;  wr_data_rom[  260]='h00000069;
    rd_cycle[  261] = 1'b0;  wr_cycle[  261] = 1'b1;  addr_rom[  261]='h00000100;  wr_data_rom[  261]='h000003c6;
    rd_cycle[  262] = 1'b1;  wr_cycle[  262] = 1'b0;  addr_rom[  262]='h000001ec;  wr_data_rom[  262]='h00000000;
    rd_cycle[  263] = 1'b0;  wr_cycle[  263] = 1'b1;  addr_rom[  263]='h00000384;  wr_data_rom[  263]='h000000a0;
    rd_cycle[  264] = 1'b1;  wr_cycle[  264] = 1'b0;  addr_rom[  264]='h000002dc;  wr_data_rom[  264]='h00000000;
    rd_cycle[  265] = 1'b0;  wr_cycle[  265] = 1'b1;  addr_rom[  265]='h00000050;  wr_data_rom[  265]='h000001ba;
    rd_cycle[  266] = 1'b0;  wr_cycle[  266] = 1'b1;  addr_rom[  266]='h00000388;  wr_data_rom[  266]='h0000007b;
    rd_cycle[  267] = 1'b0;  wr_cycle[  267] = 1'b1;  addr_rom[  267]='h000001e8;  wr_data_rom[  267]='h00000002;
    rd_cycle[  268] = 1'b1;  wr_cycle[  268] = 1'b0;  addr_rom[  268]='h00000080;  wr_data_rom[  268]='h00000000;
    rd_cycle[  269] = 1'b0;  wr_cycle[  269] = 1'b1;  addr_rom[  269]='h000002a4;  wr_data_rom[  269]='h00000106;
    rd_cycle[  270] = 1'b1;  wr_cycle[  270] = 1'b0;  addr_rom[  270]='h00000200;  wr_data_rom[  270]='h00000000;
    rd_cycle[  271] = 1'b0;  wr_cycle[  271] = 1'b1;  addr_rom[  271]='h000000bc;  wr_data_rom[  271]='h000001d7;
    rd_cycle[  272] = 1'b1;  wr_cycle[  272] = 1'b0;  addr_rom[  272]='h00000330;  wr_data_rom[  272]='h00000000;
    rd_cycle[  273] = 1'b1;  wr_cycle[  273] = 1'b0;  addr_rom[  273]='h00000144;  wr_data_rom[  273]='h00000000;
    rd_cycle[  274] = 1'b0;  wr_cycle[  274] = 1'b1;  addr_rom[  274]='h00000114;  wr_data_rom[  274]='h000001fe;
    rd_cycle[  275] = 1'b0;  wr_cycle[  275] = 1'b1;  addr_rom[  275]='h00000314;  wr_data_rom[  275]='h000002fd;
    rd_cycle[  276] = 1'b0;  wr_cycle[  276] = 1'b1;  addr_rom[  276]='h0000010c;  wr_data_rom[  276]='h00000319;
    rd_cycle[  277] = 1'b1;  wr_cycle[  277] = 1'b0;  addr_rom[  277]='h000002ec;  wr_data_rom[  277]='h00000000;
    rd_cycle[  278] = 1'b0;  wr_cycle[  278] = 1'b1;  addr_rom[  278]='h000000fc;  wr_data_rom[  278]='h00000171;
    rd_cycle[  279] = 1'b1;  wr_cycle[  279] = 1'b0;  addr_rom[  279]='h00000250;  wr_data_rom[  279]='h00000000;
    rd_cycle[  280] = 1'b0;  wr_cycle[  280] = 1'b1;  addr_rom[  280]='h0000020c;  wr_data_rom[  280]='h0000010b;
    rd_cycle[  281] = 1'b1;  wr_cycle[  281] = 1'b0;  addr_rom[  281]='h000000f8;  wr_data_rom[  281]='h00000000;
    rd_cycle[  282] = 1'b0;  wr_cycle[  282] = 1'b1;  addr_rom[  282]='h000000b4;  wr_data_rom[  282]='h000001d5;
    rd_cycle[  283] = 1'b1;  wr_cycle[  283] = 1'b0;  addr_rom[  283]='h000003a8;  wr_data_rom[  283]='h00000000;
    rd_cycle[  284] = 1'b1;  wr_cycle[  284] = 1'b0;  addr_rom[  284]='h00000080;  wr_data_rom[  284]='h00000000;
    rd_cycle[  285] = 1'b0;  wr_cycle[  285] = 1'b1;  addr_rom[  285]='h0000028c;  wr_data_rom[  285]='h000002c3;
    rd_cycle[  286] = 1'b0;  wr_cycle[  286] = 1'b1;  addr_rom[  286]='h000002c0;  wr_data_rom[  286]='h000001cc;
    rd_cycle[  287] = 1'b0;  wr_cycle[  287] = 1'b1;  addr_rom[  287]='h000000b4;  wr_data_rom[  287]='h0000025e;
    rd_cycle[  288] = 1'b0;  wr_cycle[  288] = 1'b1;  addr_rom[  288]='h00000370;  wr_data_rom[  288]='h000002d1;
    rd_cycle[  289] = 1'b0;  wr_cycle[  289] = 1'b1;  addr_rom[  289]='h00000074;  wr_data_rom[  289]='h000000e1;
    rd_cycle[  290] = 1'b1;  wr_cycle[  290] = 1'b0;  addr_rom[  290]='h00000010;  wr_data_rom[  290]='h00000000;
    rd_cycle[  291] = 1'b1;  wr_cycle[  291] = 1'b0;  addr_rom[  291]='h0000026c;  wr_data_rom[  291]='h00000000;
    rd_cycle[  292] = 1'b1;  wr_cycle[  292] = 1'b0;  addr_rom[  292]='h00000258;  wr_data_rom[  292]='h00000000;
    rd_cycle[  293] = 1'b0;  wr_cycle[  293] = 1'b1;  addr_rom[  293]='h000003f0;  wr_data_rom[  293]='h0000039f;
    rd_cycle[  294] = 1'b0;  wr_cycle[  294] = 1'b1;  addr_rom[  294]='h000000f0;  wr_data_rom[  294]='h000000b4;
    rd_cycle[  295] = 1'b1;  wr_cycle[  295] = 1'b0;  addr_rom[  295]='h00000364;  wr_data_rom[  295]='h00000000;
    rd_cycle[  296] = 1'b0;  wr_cycle[  296] = 1'b1;  addr_rom[  296]='h00000074;  wr_data_rom[  296]='h00000160;
    rd_cycle[  297] = 1'b1;  wr_cycle[  297] = 1'b0;  addr_rom[  297]='h000003e0;  wr_data_rom[  297]='h00000000;
    rd_cycle[  298] = 1'b0;  wr_cycle[  298] = 1'b1;  addr_rom[  298]='h000000a4;  wr_data_rom[  298]='h00000191;
    rd_cycle[  299] = 1'b0;  wr_cycle[  299] = 1'b1;  addr_rom[  299]='h00000018;  wr_data_rom[  299]='h00000230;
    rd_cycle[  300] = 1'b0;  wr_cycle[  300] = 1'b1;  addr_rom[  300]='h000003b8;  wr_data_rom[  300]='h00000309;
    rd_cycle[  301] = 1'b1;  wr_cycle[  301] = 1'b0;  addr_rom[  301]='h0000033c;  wr_data_rom[  301]='h00000000;
    rd_cycle[  302] = 1'b1;  wr_cycle[  302] = 1'b0;  addr_rom[  302]='h00000150;  wr_data_rom[  302]='h00000000;
    rd_cycle[  303] = 1'b1;  wr_cycle[  303] = 1'b0;  addr_rom[  303]='h00000204;  wr_data_rom[  303]='h00000000;
    rd_cycle[  304] = 1'b1;  wr_cycle[  304] = 1'b0;  addr_rom[  304]='h00000388;  wr_data_rom[  304]='h00000000;
    rd_cycle[  305] = 1'b1;  wr_cycle[  305] = 1'b0;  addr_rom[  305]='h00000274;  wr_data_rom[  305]='h00000000;
    rd_cycle[  306] = 1'b0;  wr_cycle[  306] = 1'b1;  addr_rom[  306]='h00000360;  wr_data_rom[  306]='h00000067;
    rd_cycle[  307] = 1'b1;  wr_cycle[  307] = 1'b0;  addr_rom[  307]='h00000000;  wr_data_rom[  307]='h00000000;
    rd_cycle[  308] = 1'b1;  wr_cycle[  308] = 1'b0;  addr_rom[  308]='h00000234;  wr_data_rom[  308]='h00000000;
    rd_cycle[  309] = 1'b1;  wr_cycle[  309] = 1'b0;  addr_rom[  309]='h00000124;  wr_data_rom[  309]='h00000000;
    rd_cycle[  310] = 1'b1;  wr_cycle[  310] = 1'b0;  addr_rom[  310]='h000001b4;  wr_data_rom[  310]='h00000000;
    rd_cycle[  311] = 1'b0;  wr_cycle[  311] = 1'b1;  addr_rom[  311]='h00000174;  wr_data_rom[  311]='h000002b0;
    rd_cycle[  312] = 1'b1;  wr_cycle[  312] = 1'b0;  addr_rom[  312]='h00000160;  wr_data_rom[  312]='h00000000;
    rd_cycle[  313] = 1'b0;  wr_cycle[  313] = 1'b1;  addr_rom[  313]='h0000039c;  wr_data_rom[  313]='h000002e9;
    rd_cycle[  314] = 1'b1;  wr_cycle[  314] = 1'b0;  addr_rom[  314]='h00000280;  wr_data_rom[  314]='h00000000;
    rd_cycle[  315] = 1'b0;  wr_cycle[  315] = 1'b1;  addr_rom[  315]='h0000032c;  wr_data_rom[  315]='h000000d8;
    rd_cycle[  316] = 1'b1;  wr_cycle[  316] = 1'b0;  addr_rom[  316]='h0000001c;  wr_data_rom[  316]='h00000000;
    rd_cycle[  317] = 1'b1;  wr_cycle[  317] = 1'b0;  addr_rom[  317]='h0000037c;  wr_data_rom[  317]='h00000000;
    rd_cycle[  318] = 1'b0;  wr_cycle[  318] = 1'b1;  addr_rom[  318]='h00000340;  wr_data_rom[  318]='h00000344;
    rd_cycle[  319] = 1'b1;  wr_cycle[  319] = 1'b0;  addr_rom[  319]='h000003c0;  wr_data_rom[  319]='h00000000;
    rd_cycle[  320] = 1'b0;  wr_cycle[  320] = 1'b1;  addr_rom[  320]='h00000090;  wr_data_rom[  320]='h000000f3;
    rd_cycle[  321] = 1'b0;  wr_cycle[  321] = 1'b1;  addr_rom[  321]='h00000074;  wr_data_rom[  321]='h0000031e;
    rd_cycle[  322] = 1'b0;  wr_cycle[  322] = 1'b1;  addr_rom[  322]='h00000120;  wr_data_rom[  322]='h000000f1;
    rd_cycle[  323] = 1'b0;  wr_cycle[  323] = 1'b1;  addr_rom[  323]='h00000388;  wr_data_rom[  323]='h00000400;
    rd_cycle[  324] = 1'b0;  wr_cycle[  324] = 1'b1;  addr_rom[  324]='h0000014c;  wr_data_rom[  324]='h000003cc;
    rd_cycle[  325] = 1'b1;  wr_cycle[  325] = 1'b0;  addr_rom[  325]='h00000394;  wr_data_rom[  325]='h00000000;
    rd_cycle[  326] = 1'b0;  wr_cycle[  326] = 1'b1;  addr_rom[  326]='h00000268;  wr_data_rom[  326]='h00000239;
    rd_cycle[  327] = 1'b0;  wr_cycle[  327] = 1'b1;  addr_rom[  327]='h00000020;  wr_data_rom[  327]='h000000ee;
    rd_cycle[  328] = 1'b1;  wr_cycle[  328] = 1'b0;  addr_rom[  328]='h000003ac;  wr_data_rom[  328]='h00000000;
    rd_cycle[  329] = 1'b1;  wr_cycle[  329] = 1'b0;  addr_rom[  329]='h0000027c;  wr_data_rom[  329]='h00000000;
    rd_cycle[  330] = 1'b1;  wr_cycle[  330] = 1'b0;  addr_rom[  330]='h00000098;  wr_data_rom[  330]='h00000000;
    rd_cycle[  331] = 1'b0;  wr_cycle[  331] = 1'b1;  addr_rom[  331]='h0000016c;  wr_data_rom[  331]='h0000032f;
    rd_cycle[  332] = 1'b0;  wr_cycle[  332] = 1'b1;  addr_rom[  332]='h00000078;  wr_data_rom[  332]='h00000028;
    rd_cycle[  333] = 1'b0;  wr_cycle[  333] = 1'b1;  addr_rom[  333]='h000001ec;  wr_data_rom[  333]='h000001fd;
    rd_cycle[  334] = 1'b0;  wr_cycle[  334] = 1'b1;  addr_rom[  334]='h0000003c;  wr_data_rom[  334]='h0000035f;
    rd_cycle[  335] = 1'b1;  wr_cycle[  335] = 1'b0;  addr_rom[  335]='h00000374;  wr_data_rom[  335]='h00000000;
    rd_cycle[  336] = 1'b1;  wr_cycle[  336] = 1'b0;  addr_rom[  336]='h000001bc;  wr_data_rom[  336]='h00000000;
    rd_cycle[  337] = 1'b0;  wr_cycle[  337] = 1'b1;  addr_rom[  337]='h000003d8;  wr_data_rom[  337]='h00000114;
    rd_cycle[  338] = 1'b0;  wr_cycle[  338] = 1'b1;  addr_rom[  338]='h00000324;  wr_data_rom[  338]='h00000268;
    rd_cycle[  339] = 1'b1;  wr_cycle[  339] = 1'b0;  addr_rom[  339]='h0000018c;  wr_data_rom[  339]='h00000000;
    rd_cycle[  340] = 1'b1;  wr_cycle[  340] = 1'b0;  addr_rom[  340]='h0000007c;  wr_data_rom[  340]='h00000000;
    rd_cycle[  341] = 1'b1;  wr_cycle[  341] = 1'b0;  addr_rom[  341]='h00000204;  wr_data_rom[  341]='h00000000;
    rd_cycle[  342] = 1'b1;  wr_cycle[  342] = 1'b0;  addr_rom[  342]='h00000114;  wr_data_rom[  342]='h00000000;
    rd_cycle[  343] = 1'b0;  wr_cycle[  343] = 1'b1;  addr_rom[  343]='h00000090;  wr_data_rom[  343]='h000000bb;
    rd_cycle[  344] = 1'b1;  wr_cycle[  344] = 1'b0;  addr_rom[  344]='h0000007c;  wr_data_rom[  344]='h00000000;
    rd_cycle[  345] = 1'b1;  wr_cycle[  345] = 1'b0;  addr_rom[  345]='h00000034;  wr_data_rom[  345]='h00000000;
    rd_cycle[  346] = 1'b1;  wr_cycle[  346] = 1'b0;  addr_rom[  346]='h00000174;  wr_data_rom[  346]='h00000000;
    rd_cycle[  347] = 1'b1;  wr_cycle[  347] = 1'b0;  addr_rom[  347]='h00000264;  wr_data_rom[  347]='h00000000;
    rd_cycle[  348] = 1'b1;  wr_cycle[  348] = 1'b0;  addr_rom[  348]='h00000134;  wr_data_rom[  348]='h00000000;
    rd_cycle[  349] = 1'b0;  wr_cycle[  349] = 1'b1;  addr_rom[  349]='h00000364;  wr_data_rom[  349]='h00000229;
    rd_cycle[  350] = 1'b0;  wr_cycle[  350] = 1'b1;  addr_rom[  350]='h000000ec;  wr_data_rom[  350]='h000002ff;
    rd_cycle[  351] = 1'b1;  wr_cycle[  351] = 1'b0;  addr_rom[  351]='h000002a8;  wr_data_rom[  351]='h00000000;
    rd_cycle[  352] = 1'b1;  wr_cycle[  352] = 1'b0;  addr_rom[  352]='h00000330;  wr_data_rom[  352]='h00000000;
    rd_cycle[  353] = 1'b0;  wr_cycle[  353] = 1'b1;  addr_rom[  353]='h000001dc;  wr_data_rom[  353]='h000003b8;
    rd_cycle[  354] = 1'b1;  wr_cycle[  354] = 1'b0;  addr_rom[  354]='h000002fc;  wr_data_rom[  354]='h00000000;
    rd_cycle[  355] = 1'b1;  wr_cycle[  355] = 1'b0;  addr_rom[  355]='h00000130;  wr_data_rom[  355]='h00000000;
    rd_cycle[  356] = 1'b1;  wr_cycle[  356] = 1'b0;  addr_rom[  356]='h000001d0;  wr_data_rom[  356]='h00000000;
    rd_cycle[  357] = 1'b0;  wr_cycle[  357] = 1'b1;  addr_rom[  357]='h0000010c;  wr_data_rom[  357]='h0000014a;
    rd_cycle[  358] = 1'b1;  wr_cycle[  358] = 1'b0;  addr_rom[  358]='h00000078;  wr_data_rom[  358]='h00000000;
    rd_cycle[  359] = 1'b1;  wr_cycle[  359] = 1'b0;  addr_rom[  359]='h0000031c;  wr_data_rom[  359]='h00000000;
    rd_cycle[  360] = 1'b1;  wr_cycle[  360] = 1'b0;  addr_rom[  360]='h00000284;  wr_data_rom[  360]='h00000000;
    rd_cycle[  361] = 1'b1;  wr_cycle[  361] = 1'b0;  addr_rom[  361]='h000002c4;  wr_data_rom[  361]='h00000000;
    rd_cycle[  362] = 1'b0;  wr_cycle[  362] = 1'b1;  addr_rom[  362]='h0000013c;  wr_data_rom[  362]='h00000224;
    rd_cycle[  363] = 1'b1;  wr_cycle[  363] = 1'b0;  addr_rom[  363]='h000003bc;  wr_data_rom[  363]='h00000000;
    rd_cycle[  364] = 1'b1;  wr_cycle[  364] = 1'b0;  addr_rom[  364]='h00000304;  wr_data_rom[  364]='h00000000;
    rd_cycle[  365] = 1'b1;  wr_cycle[  365] = 1'b0;  addr_rom[  365]='h000001c0;  wr_data_rom[  365]='h00000000;
    rd_cycle[  366] = 1'b1;  wr_cycle[  366] = 1'b0;  addr_rom[  366]='h00000268;  wr_data_rom[  366]='h00000000;
    rd_cycle[  367] = 1'b1;  wr_cycle[  367] = 1'b0;  addr_rom[  367]='h00000198;  wr_data_rom[  367]='h00000000;
    rd_cycle[  368] = 1'b0;  wr_cycle[  368] = 1'b1;  addr_rom[  368]='h00000048;  wr_data_rom[  368]='h00000335;
    rd_cycle[  369] = 1'b0;  wr_cycle[  369] = 1'b1;  addr_rom[  369]='h000002a8;  wr_data_rom[  369]='h000000e5;
    rd_cycle[  370] = 1'b0;  wr_cycle[  370] = 1'b1;  addr_rom[  370]='h000002b4;  wr_data_rom[  370]='h00000339;
    rd_cycle[  371] = 1'b1;  wr_cycle[  371] = 1'b0;  addr_rom[  371]='h00000130;  wr_data_rom[  371]='h00000000;
    rd_cycle[  372] = 1'b1;  wr_cycle[  372] = 1'b0;  addr_rom[  372]='h000000a4;  wr_data_rom[  372]='h00000000;
    rd_cycle[  373] = 1'b1;  wr_cycle[  373] = 1'b0;  addr_rom[  373]='h00000330;  wr_data_rom[  373]='h00000000;
    rd_cycle[  374] = 1'b1;  wr_cycle[  374] = 1'b0;  addr_rom[  374]='h0000004c;  wr_data_rom[  374]='h00000000;
    rd_cycle[  375] = 1'b1;  wr_cycle[  375] = 1'b0;  addr_rom[  375]='h00000220;  wr_data_rom[  375]='h00000000;
    rd_cycle[  376] = 1'b0;  wr_cycle[  376] = 1'b1;  addr_rom[  376]='h00000144;  wr_data_rom[  376]='h000002f3;
    rd_cycle[  377] = 1'b0;  wr_cycle[  377] = 1'b1;  addr_rom[  377]='h00000248;  wr_data_rom[  377]='h00000062;
    rd_cycle[  378] = 1'b0;  wr_cycle[  378] = 1'b1;  addr_rom[  378]='h000002c0;  wr_data_rom[  378]='h00000224;
    rd_cycle[  379] = 1'b1;  wr_cycle[  379] = 1'b0;  addr_rom[  379]='h000000e0;  wr_data_rom[  379]='h00000000;
    rd_cycle[  380] = 1'b1;  wr_cycle[  380] = 1'b0;  addr_rom[  380]='h000002c0;  wr_data_rom[  380]='h00000000;
    rd_cycle[  381] = 1'b1;  wr_cycle[  381] = 1'b0;  addr_rom[  381]='h00000190;  wr_data_rom[  381]='h00000000;
    rd_cycle[  382] = 1'b0;  wr_cycle[  382] = 1'b1;  addr_rom[  382]='h000000f4;  wr_data_rom[  382]='h00000304;
    rd_cycle[  383] = 1'b0;  wr_cycle[  383] = 1'b1;  addr_rom[  383]='h00000220;  wr_data_rom[  383]='h000000ca;
    rd_cycle[  384] = 1'b0;  wr_cycle[  384] = 1'b1;  addr_rom[  384]='h000001d4;  wr_data_rom[  384]='h00000345;
    rd_cycle[  385] = 1'b1;  wr_cycle[  385] = 1'b0;  addr_rom[  385]='h000001b0;  wr_data_rom[  385]='h00000000;
    rd_cycle[  386] = 1'b1;  wr_cycle[  386] = 1'b0;  addr_rom[  386]='h00000310;  wr_data_rom[  386]='h00000000;
    rd_cycle[  387] = 1'b0;  wr_cycle[  387] = 1'b1;  addr_rom[  387]='h0000007c;  wr_data_rom[  387]='h0000004a;
    rd_cycle[  388] = 1'b1;  wr_cycle[  388] = 1'b0;  addr_rom[  388]='h00000398;  wr_data_rom[  388]='h00000000;
    rd_cycle[  389] = 1'b0;  wr_cycle[  389] = 1'b1;  addr_rom[  389]='h00000000;  wr_data_rom[  389]='h000001a9;
    rd_cycle[  390] = 1'b0;  wr_cycle[  390] = 1'b1;  addr_rom[  390]='h000003bc;  wr_data_rom[  390]='h000001ca;
    rd_cycle[  391] = 1'b0;  wr_cycle[  391] = 1'b1;  addr_rom[  391]='h000003b8;  wr_data_rom[  391]='h000001a7;
    rd_cycle[  392] = 1'b0;  wr_cycle[  392] = 1'b1;  addr_rom[  392]='h00000358;  wr_data_rom[  392]='h00000236;
    rd_cycle[  393] = 1'b0;  wr_cycle[  393] = 1'b1;  addr_rom[  393]='h000001e0;  wr_data_rom[  393]='h000002f1;
    rd_cycle[  394] = 1'b0;  wr_cycle[  394] = 1'b1;  addr_rom[  394]='h0000031c;  wr_data_rom[  394]='h000003ee;
    rd_cycle[  395] = 1'b0;  wr_cycle[  395] = 1'b1;  addr_rom[  395]='h0000030c;  wr_data_rom[  395]='h0000008e;
    rd_cycle[  396] = 1'b0;  wr_cycle[  396] = 1'b1;  addr_rom[  396]='h000001e0;  wr_data_rom[  396]='h0000007e;
    rd_cycle[  397] = 1'b1;  wr_cycle[  397] = 1'b0;  addr_rom[  397]='h0000007c;  wr_data_rom[  397]='h00000000;
    rd_cycle[  398] = 1'b1;  wr_cycle[  398] = 1'b0;  addr_rom[  398]='h00000388;  wr_data_rom[  398]='h00000000;
    rd_cycle[  399] = 1'b1;  wr_cycle[  399] = 1'b0;  addr_rom[  399]='h00000128;  wr_data_rom[  399]='h00000000;
    rd_cycle[  400] = 1'b1;  wr_cycle[  400] = 1'b0;  addr_rom[  400]='h00000354;  wr_data_rom[  400]='h00000000;
    rd_cycle[  401] = 1'b1;  wr_cycle[  401] = 1'b0;  addr_rom[  401]='h000002e8;  wr_data_rom[  401]='h00000000;
    rd_cycle[  402] = 1'b1;  wr_cycle[  402] = 1'b0;  addr_rom[  402]='h00000224;  wr_data_rom[  402]='h00000000;
    rd_cycle[  403] = 1'b1;  wr_cycle[  403] = 1'b0;  addr_rom[  403]='h000002a4;  wr_data_rom[  403]='h00000000;
    rd_cycle[  404] = 1'b1;  wr_cycle[  404] = 1'b0;  addr_rom[  404]='h00000184;  wr_data_rom[  404]='h00000000;
    rd_cycle[  405] = 1'b0;  wr_cycle[  405] = 1'b1;  addr_rom[  405]='h000002d8;  wr_data_rom[  405]='h00000162;
    rd_cycle[  406] = 1'b1;  wr_cycle[  406] = 1'b0;  addr_rom[  406]='h00000220;  wr_data_rom[  406]='h00000000;
    rd_cycle[  407] = 1'b1;  wr_cycle[  407] = 1'b0;  addr_rom[  407]='h00000294;  wr_data_rom[  407]='h00000000;
    rd_cycle[  408] = 1'b0;  wr_cycle[  408] = 1'b1;  addr_rom[  408]='h00000358;  wr_data_rom[  408]='h000001f0;
    rd_cycle[  409] = 1'b1;  wr_cycle[  409] = 1'b0;  addr_rom[  409]='h0000022c;  wr_data_rom[  409]='h00000000;
    rd_cycle[  410] = 1'b1;  wr_cycle[  410] = 1'b0;  addr_rom[  410]='h00000290;  wr_data_rom[  410]='h00000000;
    rd_cycle[  411] = 1'b0;  wr_cycle[  411] = 1'b1;  addr_rom[  411]='h0000007c;  wr_data_rom[  411]='h00000034;
    rd_cycle[  412] = 1'b1;  wr_cycle[  412] = 1'b0;  addr_rom[  412]='h000001a8;  wr_data_rom[  412]='h00000000;
    rd_cycle[  413] = 1'b0;  wr_cycle[  413] = 1'b1;  addr_rom[  413]='h000003d0;  wr_data_rom[  413]='h0000018c;
    rd_cycle[  414] = 1'b0;  wr_cycle[  414] = 1'b1;  addr_rom[  414]='h00000024;  wr_data_rom[  414]='h00000280;
    rd_cycle[  415] = 1'b1;  wr_cycle[  415] = 1'b0;  addr_rom[  415]='h00000024;  wr_data_rom[  415]='h00000000;
    rd_cycle[  416] = 1'b0;  wr_cycle[  416] = 1'b1;  addr_rom[  416]='h00000254;  wr_data_rom[  416]='h0000034b;
    rd_cycle[  417] = 1'b1;  wr_cycle[  417] = 1'b0;  addr_rom[  417]='h0000007c;  wr_data_rom[  417]='h00000000;
    rd_cycle[  418] = 1'b0;  wr_cycle[  418] = 1'b1;  addr_rom[  418]='h000003b4;  wr_data_rom[  418]='h00000226;
    rd_cycle[  419] = 1'b1;  wr_cycle[  419] = 1'b0;  addr_rom[  419]='h00000214;  wr_data_rom[  419]='h00000000;
    rd_cycle[  420] = 1'b0;  wr_cycle[  420] = 1'b1;  addr_rom[  420]='h0000034c;  wr_data_rom[  420]='h000002f9;
    rd_cycle[  421] = 1'b1;  wr_cycle[  421] = 1'b0;  addr_rom[  421]='h0000007c;  wr_data_rom[  421]='h00000000;
    rd_cycle[  422] = 1'b1;  wr_cycle[  422] = 1'b0;  addr_rom[  422]='h000002a0;  wr_data_rom[  422]='h00000000;
    rd_cycle[  423] = 1'b0;  wr_cycle[  423] = 1'b1;  addr_rom[  423]='h000002d8;  wr_data_rom[  423]='h000001fe;
    rd_cycle[  424] = 1'b1;  wr_cycle[  424] = 1'b0;  addr_rom[  424]='h00000164;  wr_data_rom[  424]='h00000000;
    rd_cycle[  425] = 1'b1;  wr_cycle[  425] = 1'b0;  addr_rom[  425]='h000003e8;  wr_data_rom[  425]='h00000000;
    rd_cycle[  426] = 1'b1;  wr_cycle[  426] = 1'b0;  addr_rom[  426]='h00000240;  wr_data_rom[  426]='h00000000;
    rd_cycle[  427] = 1'b1;  wr_cycle[  427] = 1'b0;  addr_rom[  427]='h00000368;  wr_data_rom[  427]='h00000000;
    rd_cycle[  428] = 1'b1;  wr_cycle[  428] = 1'b0;  addr_rom[  428]='h000002cc;  wr_data_rom[  428]='h00000000;
    rd_cycle[  429] = 1'b0;  wr_cycle[  429] = 1'b1;  addr_rom[  429]='h0000036c;  wr_data_rom[  429]='h000002fb;
    rd_cycle[  430] = 1'b0;  wr_cycle[  430] = 1'b1;  addr_rom[  430]='h000000a8;  wr_data_rom[  430]='h00000130;
    rd_cycle[  431] = 1'b0;  wr_cycle[  431] = 1'b1;  addr_rom[  431]='h000000f0;  wr_data_rom[  431]='h000002d4;
    rd_cycle[  432] = 1'b0;  wr_cycle[  432] = 1'b1;  addr_rom[  432]='h00000178;  wr_data_rom[  432]='h0000001c;
    rd_cycle[  433] = 1'b1;  wr_cycle[  433] = 1'b0;  addr_rom[  433]='h000002d0;  wr_data_rom[  433]='h00000000;
    rd_cycle[  434] = 1'b0;  wr_cycle[  434] = 1'b1;  addr_rom[  434]='h000003a4;  wr_data_rom[  434]='h0000014c;
    rd_cycle[  435] = 1'b1;  wr_cycle[  435] = 1'b0;  addr_rom[  435]='h000001d8;  wr_data_rom[  435]='h00000000;
    rd_cycle[  436] = 1'b1;  wr_cycle[  436] = 1'b0;  addr_rom[  436]='h000000f8;  wr_data_rom[  436]='h00000000;
    rd_cycle[  437] = 1'b0;  wr_cycle[  437] = 1'b1;  addr_rom[  437]='h0000031c;  wr_data_rom[  437]='h00000178;
    rd_cycle[  438] = 1'b1;  wr_cycle[  438] = 1'b0;  addr_rom[  438]='h00000378;  wr_data_rom[  438]='h00000000;
    rd_cycle[  439] = 1'b1;  wr_cycle[  439] = 1'b0;  addr_rom[  439]='h000000e0;  wr_data_rom[  439]='h00000000;
    rd_cycle[  440] = 1'b1;  wr_cycle[  440] = 1'b0;  addr_rom[  440]='h00000124;  wr_data_rom[  440]='h00000000;
    rd_cycle[  441] = 1'b1;  wr_cycle[  441] = 1'b0;  addr_rom[  441]='h000002f4;  wr_data_rom[  441]='h00000000;
    rd_cycle[  442] = 1'b1;  wr_cycle[  442] = 1'b0;  addr_rom[  442]='h0000036c;  wr_data_rom[  442]='h00000000;
    rd_cycle[  443] = 1'b1;  wr_cycle[  443] = 1'b0;  addr_rom[  443]='h00000288;  wr_data_rom[  443]='h00000000;
    rd_cycle[  444] = 1'b0;  wr_cycle[  444] = 1'b1;  addr_rom[  444]='h00000368;  wr_data_rom[  444]='h000001f1;
    rd_cycle[  445] = 1'b1;  wr_cycle[  445] = 1'b0;  addr_rom[  445]='h00000370;  wr_data_rom[  445]='h00000000;
    rd_cycle[  446] = 1'b1;  wr_cycle[  446] = 1'b0;  addr_rom[  446]='h000000a0;  wr_data_rom[  446]='h00000000;
    rd_cycle[  447] = 1'b1;  wr_cycle[  447] = 1'b0;  addr_rom[  447]='h000003d4;  wr_data_rom[  447]='h00000000;
    rd_cycle[  448] = 1'b0;  wr_cycle[  448] = 1'b1;  addr_rom[  448]='h00000218;  wr_data_rom[  448]='h00000216;
    rd_cycle[  449] = 1'b0;  wr_cycle[  449] = 1'b1;  addr_rom[  449]='h0000005c;  wr_data_rom[  449]='h00000025;
    rd_cycle[  450] = 1'b1;  wr_cycle[  450] = 1'b0;  addr_rom[  450]='h000001c0;  wr_data_rom[  450]='h00000000;
    rd_cycle[  451] = 1'b0;  wr_cycle[  451] = 1'b1;  addr_rom[  451]='h00000010;  wr_data_rom[  451]='h0000034f;
    rd_cycle[  452] = 1'b0;  wr_cycle[  452] = 1'b1;  addr_rom[  452]='h0000032c;  wr_data_rom[  452]='h0000025a;
    rd_cycle[  453] = 1'b0;  wr_cycle[  453] = 1'b1;  addr_rom[  453]='h00000250;  wr_data_rom[  453]='h00000249;
    rd_cycle[  454] = 1'b1;  wr_cycle[  454] = 1'b0;  addr_rom[  454]='h000003a4;  wr_data_rom[  454]='h00000000;
    rd_cycle[  455] = 1'b1;  wr_cycle[  455] = 1'b0;  addr_rom[  455]='h000000b0;  wr_data_rom[  455]='h00000000;
    rd_cycle[  456] = 1'b1;  wr_cycle[  456] = 1'b0;  addr_rom[  456]='h000003c0;  wr_data_rom[  456]='h00000000;
    rd_cycle[  457] = 1'b1;  wr_cycle[  457] = 1'b0;  addr_rom[  457]='h0000021c;  wr_data_rom[  457]='h00000000;
    rd_cycle[  458] = 1'b0;  wr_cycle[  458] = 1'b1;  addr_rom[  458]='h00000110;  wr_data_rom[  458]='h00000259;
    rd_cycle[  459] = 1'b0;  wr_cycle[  459] = 1'b1;  addr_rom[  459]='h00000340;  wr_data_rom[  459]='h0000031f;
    rd_cycle[  460] = 1'b0;  wr_cycle[  460] = 1'b1;  addr_rom[  460]='h00000120;  wr_data_rom[  460]='h00000314;
    rd_cycle[  461] = 1'b0;  wr_cycle[  461] = 1'b1;  addr_rom[  461]='h000000c8;  wr_data_rom[  461]='h000001ef;
    rd_cycle[  462] = 1'b1;  wr_cycle[  462] = 1'b0;  addr_rom[  462]='h000003ec;  wr_data_rom[  462]='h00000000;
    rd_cycle[  463] = 1'b1;  wr_cycle[  463] = 1'b0;  addr_rom[  463]='h00000060;  wr_data_rom[  463]='h00000000;
    rd_cycle[  464] = 1'b0;  wr_cycle[  464] = 1'b1;  addr_rom[  464]='h00000144;  wr_data_rom[  464]='h00000327;
    rd_cycle[  465] = 1'b1;  wr_cycle[  465] = 1'b0;  addr_rom[  465]='h000000b8;  wr_data_rom[  465]='h00000000;
    rd_cycle[  466] = 1'b1;  wr_cycle[  466] = 1'b0;  addr_rom[  466]='h00000108;  wr_data_rom[  466]='h00000000;
    rd_cycle[  467] = 1'b1;  wr_cycle[  467] = 1'b0;  addr_rom[  467]='h0000020c;  wr_data_rom[  467]='h00000000;
    rd_cycle[  468] = 1'b0;  wr_cycle[  468] = 1'b1;  addr_rom[  468]='h000001f4;  wr_data_rom[  468]='h000000b2;
    rd_cycle[  469] = 1'b0;  wr_cycle[  469] = 1'b1;  addr_rom[  469]='h000000e8;  wr_data_rom[  469]='h00000364;
    rd_cycle[  470] = 1'b1;  wr_cycle[  470] = 1'b0;  addr_rom[  470]='h00000134;  wr_data_rom[  470]='h00000000;
    rd_cycle[  471] = 1'b1;  wr_cycle[  471] = 1'b0;  addr_rom[  471]='h000001c8;  wr_data_rom[  471]='h00000000;
    rd_cycle[  472] = 1'b0;  wr_cycle[  472] = 1'b1;  addr_rom[  472]='h00000098;  wr_data_rom[  472]='h0000003a;
    rd_cycle[  473] = 1'b1;  wr_cycle[  473] = 1'b0;  addr_rom[  473]='h0000034c;  wr_data_rom[  473]='h00000000;
    rd_cycle[  474] = 1'b0;  wr_cycle[  474] = 1'b1;  addr_rom[  474]='h000000b0;  wr_data_rom[  474]='h000003a3;
    rd_cycle[  475] = 1'b0;  wr_cycle[  475] = 1'b1;  addr_rom[  475]='h000001bc;  wr_data_rom[  475]='h00000070;
    rd_cycle[  476] = 1'b0;  wr_cycle[  476] = 1'b1;  addr_rom[  476]='h000000b0;  wr_data_rom[  476]='h0000028d;
    rd_cycle[  477] = 1'b0;  wr_cycle[  477] = 1'b1;  addr_rom[  477]='h00000178;  wr_data_rom[  477]='h000002a7;
    rd_cycle[  478] = 1'b0;  wr_cycle[  478] = 1'b1;  addr_rom[  478]='h000002d4;  wr_data_rom[  478]='h00000291;
    rd_cycle[  479] = 1'b0;  wr_cycle[  479] = 1'b1;  addr_rom[  479]='h000000e0;  wr_data_rom[  479]='h0000016f;
    rd_cycle[  480] = 1'b1;  wr_cycle[  480] = 1'b0;  addr_rom[  480]='h0000024c;  wr_data_rom[  480]='h00000000;
    rd_cycle[  481] = 1'b0;  wr_cycle[  481] = 1'b1;  addr_rom[  481]='h00000288;  wr_data_rom[  481]='h00000041;
    rd_cycle[  482] = 1'b0;  wr_cycle[  482] = 1'b1;  addr_rom[  482]='h000001e4;  wr_data_rom[  482]='h000001f6;
    rd_cycle[  483] = 1'b1;  wr_cycle[  483] = 1'b0;  addr_rom[  483]='h00000038;  wr_data_rom[  483]='h00000000;
    rd_cycle[  484] = 1'b1;  wr_cycle[  484] = 1'b0;  addr_rom[  484]='h000000f0;  wr_data_rom[  484]='h00000000;
    rd_cycle[  485] = 1'b1;  wr_cycle[  485] = 1'b0;  addr_rom[  485]='h00000378;  wr_data_rom[  485]='h00000000;
    rd_cycle[  486] = 1'b0;  wr_cycle[  486] = 1'b1;  addr_rom[  486]='h000002d0;  wr_data_rom[  486]='h000003ce;
    rd_cycle[  487] = 1'b1;  wr_cycle[  487] = 1'b0;  addr_rom[  487]='h00000238;  wr_data_rom[  487]='h00000000;
    rd_cycle[  488] = 1'b1;  wr_cycle[  488] = 1'b0;  addr_rom[  488]='h00000124;  wr_data_rom[  488]='h00000000;
    rd_cycle[  489] = 1'b1;  wr_cycle[  489] = 1'b0;  addr_rom[  489]='h000000b0;  wr_data_rom[  489]='h00000000;
    rd_cycle[  490] = 1'b1;  wr_cycle[  490] = 1'b0;  addr_rom[  490]='h000001d4;  wr_data_rom[  490]='h00000000;
    rd_cycle[  491] = 1'b0;  wr_cycle[  491] = 1'b1;  addr_rom[  491]='h00000138;  wr_data_rom[  491]='h000000db;
    rd_cycle[  492] = 1'b1;  wr_cycle[  492] = 1'b0;  addr_rom[  492]='h00000120;  wr_data_rom[  492]='h00000000;
    rd_cycle[  493] = 1'b1;  wr_cycle[  493] = 1'b0;  addr_rom[  493]='h00000040;  wr_data_rom[  493]='h00000000;
    rd_cycle[  494] = 1'b1;  wr_cycle[  494] = 1'b0;  addr_rom[  494]='h000003a0;  wr_data_rom[  494]='h00000000;
    rd_cycle[  495] = 1'b1;  wr_cycle[  495] = 1'b0;  addr_rom[  495]='h000000b8;  wr_data_rom[  495]='h00000000;
    rd_cycle[  496] = 1'b1;  wr_cycle[  496] = 1'b0;  addr_rom[  496]='h00000264;  wr_data_rom[  496]='h00000000;
    rd_cycle[  497] = 1'b1;  wr_cycle[  497] = 1'b0;  addr_rom[  497]='h000001f0;  wr_data_rom[  497]='h00000000;
    rd_cycle[  498] = 1'b0;  wr_cycle[  498] = 1'b1;  addr_rom[  498]='h00000154;  wr_data_rom[  498]='h0000032e;
    rd_cycle[  499] = 1'b1;  wr_cycle[  499] = 1'b0;  addr_rom[  499]='h000001b8;  wr_data_rom[  499]='h00000000;
    rd_cycle[  500] = 1'b1;  wr_cycle[  500] = 1'b0;  addr_rom[  500]='h000002bc;  wr_data_rom[  500]='h00000000;
    rd_cycle[  501] = 1'b0;  wr_cycle[  501] = 1'b1;  addr_rom[  501]='h0000012c;  wr_data_rom[  501]='h000001f5;
    rd_cycle[  502] = 1'b0;  wr_cycle[  502] = 1'b1;  addr_rom[  502]='h00000344;  wr_data_rom[  502]='h000003af;
    rd_cycle[  503] = 1'b0;  wr_cycle[  503] = 1'b1;  addr_rom[  503]='h00000330;  wr_data_rom[  503]='h000003ca;
    rd_cycle[  504] = 1'b1;  wr_cycle[  504] = 1'b0;  addr_rom[  504]='h0000025c;  wr_data_rom[  504]='h00000000;
    rd_cycle[  505] = 1'b1;  wr_cycle[  505] = 1'b0;  addr_rom[  505]='h00000368;  wr_data_rom[  505]='h00000000;
    rd_cycle[  506] = 1'b1;  wr_cycle[  506] = 1'b0;  addr_rom[  506]='h00000140;  wr_data_rom[  506]='h00000000;
    rd_cycle[  507] = 1'b1;  wr_cycle[  507] = 1'b0;  addr_rom[  507]='h0000004c;  wr_data_rom[  507]='h00000000;
    rd_cycle[  508] = 1'b1;  wr_cycle[  508] = 1'b0;  addr_rom[  508]='h00000098;  wr_data_rom[  508]='h00000000;
    rd_cycle[  509] = 1'b1;  wr_cycle[  509] = 1'b0;  addr_rom[  509]='h0000007c;  wr_data_rom[  509]='h00000000;
    rd_cycle[  510] = 1'b1;  wr_cycle[  510] = 1'b0;  addr_rom[  510]='h00000198;  wr_data_rom[  510]='h00000000;
    rd_cycle[  511] = 1'b0;  wr_cycle[  511] = 1'b1;  addr_rom[  511]='h000000f0;  wr_data_rom[  511]='h000000d1;
    rd_cycle[  512] = 1'b0;  wr_cycle[  512] = 1'b1;  addr_rom[  512]='h00000040;  wr_data_rom[  512]='h00000178;
    rd_cycle[  513] = 1'b1;  wr_cycle[  513] = 1'b0;  addr_rom[  513]='h00000260;  wr_data_rom[  513]='h00000000;
    rd_cycle[  514] = 1'b1;  wr_cycle[  514] = 1'b0;  addr_rom[  514]='h000002b8;  wr_data_rom[  514]='h00000000;
    rd_cycle[  515] = 1'b1;  wr_cycle[  515] = 1'b0;  addr_rom[  515]='h0000017c;  wr_data_rom[  515]='h00000000;
    rd_cycle[  516] = 1'b0;  wr_cycle[  516] = 1'b1;  addr_rom[  516]='h000002e0;  wr_data_rom[  516]='h0000010c;
    rd_cycle[  517] = 1'b0;  wr_cycle[  517] = 1'b1;  addr_rom[  517]='h0000007c;  wr_data_rom[  517]='h000000eb;
    rd_cycle[  518] = 1'b0;  wr_cycle[  518] = 1'b1;  addr_rom[  518]='h00000380;  wr_data_rom[  518]='h000003cc;
    rd_cycle[  519] = 1'b1;  wr_cycle[  519] = 1'b0;  addr_rom[  519]='h0000001c;  wr_data_rom[  519]='h00000000;
    rd_cycle[  520] = 1'b1;  wr_cycle[  520] = 1'b0;  addr_rom[  520]='h00000144;  wr_data_rom[  520]='h00000000;
    rd_cycle[  521] = 1'b0;  wr_cycle[  521] = 1'b1;  addr_rom[  521]='h00000024;  wr_data_rom[  521]='h00000389;
    rd_cycle[  522] = 1'b1;  wr_cycle[  522] = 1'b0;  addr_rom[  522]='h00000328;  wr_data_rom[  522]='h00000000;
    rd_cycle[  523] = 1'b0;  wr_cycle[  523] = 1'b1;  addr_rom[  523]='h00000390;  wr_data_rom[  523]='h0000026b;
    rd_cycle[  524] = 1'b0;  wr_cycle[  524] = 1'b1;  addr_rom[  524]='h000003a4;  wr_data_rom[  524]='h0000010b;
    rd_cycle[  525] = 1'b0;  wr_cycle[  525] = 1'b1;  addr_rom[  525]='h00000148;  wr_data_rom[  525]='h00000221;
    rd_cycle[  526] = 1'b0;  wr_cycle[  526] = 1'b1;  addr_rom[  526]='h00000218;  wr_data_rom[  526]='h000000b6;
    rd_cycle[  527] = 1'b1;  wr_cycle[  527] = 1'b0;  addr_rom[  527]='h00000208;  wr_data_rom[  527]='h00000000;
    rd_cycle[  528] = 1'b1;  wr_cycle[  528] = 1'b0;  addr_rom[  528]='h000000c8;  wr_data_rom[  528]='h00000000;
    rd_cycle[  529] = 1'b0;  wr_cycle[  529] = 1'b1;  addr_rom[  529]='h0000032c;  wr_data_rom[  529]='h00000208;
    rd_cycle[  530] = 1'b1;  wr_cycle[  530] = 1'b0;  addr_rom[  530]='h00000190;  wr_data_rom[  530]='h00000000;
    rd_cycle[  531] = 1'b1;  wr_cycle[  531] = 1'b0;  addr_rom[  531]='h000002ac;  wr_data_rom[  531]='h00000000;
    rd_cycle[  532] = 1'b1;  wr_cycle[  532] = 1'b0;  addr_rom[  532]='h00000300;  wr_data_rom[  532]='h00000000;
    rd_cycle[  533] = 1'b1;  wr_cycle[  533] = 1'b0;  addr_rom[  533]='h000003f8;  wr_data_rom[  533]='h00000000;
    rd_cycle[  534] = 1'b0;  wr_cycle[  534] = 1'b1;  addr_rom[  534]='h00000250;  wr_data_rom[  534]='h00000125;
    rd_cycle[  535] = 1'b0;  wr_cycle[  535] = 1'b1;  addr_rom[  535]='h000000e0;  wr_data_rom[  535]='h00000361;
    rd_cycle[  536] = 1'b0;  wr_cycle[  536] = 1'b1;  addr_rom[  536]='h000002ac;  wr_data_rom[  536]='h0000002f;
    rd_cycle[  537] = 1'b0;  wr_cycle[  537] = 1'b1;  addr_rom[  537]='h00000084;  wr_data_rom[  537]='h00000286;
    rd_cycle[  538] = 1'b0;  wr_cycle[  538] = 1'b1;  addr_rom[  538]='h000001e0;  wr_data_rom[  538]='h000000d5;
    rd_cycle[  539] = 1'b1;  wr_cycle[  539] = 1'b0;  addr_rom[  539]='h000003f8;  wr_data_rom[  539]='h00000000;
    rd_cycle[  540] = 1'b0;  wr_cycle[  540] = 1'b1;  addr_rom[  540]='h000001a4;  wr_data_rom[  540]='h0000026a;
    rd_cycle[  541] = 1'b1;  wr_cycle[  541] = 1'b0;  addr_rom[  541]='h000003dc;  wr_data_rom[  541]='h00000000;
    rd_cycle[  542] = 1'b0;  wr_cycle[  542] = 1'b1;  addr_rom[  542]='h000000f8;  wr_data_rom[  542]='h00000138;
    rd_cycle[  543] = 1'b1;  wr_cycle[  543] = 1'b0;  addr_rom[  543]='h00000230;  wr_data_rom[  543]='h00000000;
    rd_cycle[  544] = 1'b0;  wr_cycle[  544] = 1'b1;  addr_rom[  544]='h00000210;  wr_data_rom[  544]='h000000a5;
    rd_cycle[  545] = 1'b0;  wr_cycle[  545] = 1'b1;  addr_rom[  545]='h00000324;  wr_data_rom[  545]='h000003be;
    rd_cycle[  546] = 1'b0;  wr_cycle[  546] = 1'b1;  addr_rom[  546]='h000001f4;  wr_data_rom[  546]='h00000330;
    rd_cycle[  547] = 1'b0;  wr_cycle[  547] = 1'b1;  addr_rom[  547]='h000000b0;  wr_data_rom[  547]='h00000305;
    rd_cycle[  548] = 1'b1;  wr_cycle[  548] = 1'b0;  addr_rom[  548]='h00000000;  wr_data_rom[  548]='h00000000;
    rd_cycle[  549] = 1'b0;  wr_cycle[  549] = 1'b1;  addr_rom[  549]='h00000358;  wr_data_rom[  549]='h0000026d;
    rd_cycle[  550] = 1'b0;  wr_cycle[  550] = 1'b1;  addr_rom[  550]='h00000348;  wr_data_rom[  550]='h00000221;
    rd_cycle[  551] = 1'b0;  wr_cycle[  551] = 1'b1;  addr_rom[  551]='h00000278;  wr_data_rom[  551]='h00000094;
    rd_cycle[  552] = 1'b0;  wr_cycle[  552] = 1'b1;  addr_rom[  552]='h000001cc;  wr_data_rom[  552]='h000003af;
    rd_cycle[  553] = 1'b0;  wr_cycle[  553] = 1'b1;  addr_rom[  553]='h000001cc;  wr_data_rom[  553]='h0000012a;
    rd_cycle[  554] = 1'b0;  wr_cycle[  554] = 1'b1;  addr_rom[  554]='h00000380;  wr_data_rom[  554]='h00000205;
    rd_cycle[  555] = 1'b1;  wr_cycle[  555] = 1'b0;  addr_rom[  555]='h0000038c;  wr_data_rom[  555]='h00000000;
    rd_cycle[  556] = 1'b0;  wr_cycle[  556] = 1'b1;  addr_rom[  556]='h000002c4;  wr_data_rom[  556]='h00000174;
    rd_cycle[  557] = 1'b0;  wr_cycle[  557] = 1'b1;  addr_rom[  557]='h000001cc;  wr_data_rom[  557]='h00000189;
    rd_cycle[  558] = 1'b0;  wr_cycle[  558] = 1'b1;  addr_rom[  558]='h0000000c;  wr_data_rom[  558]='h00000355;
    rd_cycle[  559] = 1'b1;  wr_cycle[  559] = 1'b0;  addr_rom[  559]='h000001cc;  wr_data_rom[  559]='h00000000;
    rd_cycle[  560] = 1'b0;  wr_cycle[  560] = 1'b1;  addr_rom[  560]='h00000294;  wr_data_rom[  560]='h000001fc;
    rd_cycle[  561] = 1'b1;  wr_cycle[  561] = 1'b0;  addr_rom[  561]='h00000330;  wr_data_rom[  561]='h00000000;
    rd_cycle[  562] = 1'b0;  wr_cycle[  562] = 1'b1;  addr_rom[  562]='h000000e8;  wr_data_rom[  562]='h000001a4;
    rd_cycle[  563] = 1'b1;  wr_cycle[  563] = 1'b0;  addr_rom[  563]='h000002cc;  wr_data_rom[  563]='h00000000;
    rd_cycle[  564] = 1'b1;  wr_cycle[  564] = 1'b0;  addr_rom[  564]='h000001f8;  wr_data_rom[  564]='h00000000;
    rd_cycle[  565] = 1'b1;  wr_cycle[  565] = 1'b0;  addr_rom[  565]='h00000064;  wr_data_rom[  565]='h00000000;
    rd_cycle[  566] = 1'b1;  wr_cycle[  566] = 1'b0;  addr_rom[  566]='h000001fc;  wr_data_rom[  566]='h00000000;
    rd_cycle[  567] = 1'b0;  wr_cycle[  567] = 1'b1;  addr_rom[  567]='h000003e8;  wr_data_rom[  567]='h00000396;
    rd_cycle[  568] = 1'b0;  wr_cycle[  568] = 1'b1;  addr_rom[  568]='h00000318;  wr_data_rom[  568]='h00000307;
    rd_cycle[  569] = 1'b1;  wr_cycle[  569] = 1'b0;  addr_rom[  569]='h00000160;  wr_data_rom[  569]='h00000000;
    rd_cycle[  570] = 1'b0;  wr_cycle[  570] = 1'b1;  addr_rom[  570]='h0000039c;  wr_data_rom[  570]='h000003be;
    rd_cycle[  571] = 1'b1;  wr_cycle[  571] = 1'b0;  addr_rom[  571]='h000001d4;  wr_data_rom[  571]='h00000000;
    rd_cycle[  572] = 1'b1;  wr_cycle[  572] = 1'b0;  addr_rom[  572]='h00000254;  wr_data_rom[  572]='h00000000;
    rd_cycle[  573] = 1'b0;  wr_cycle[  573] = 1'b1;  addr_rom[  573]='h000002b4;  wr_data_rom[  573]='h00000004;
    rd_cycle[  574] = 1'b1;  wr_cycle[  574] = 1'b0;  addr_rom[  574]='h00000040;  wr_data_rom[  574]='h00000000;
    rd_cycle[  575] = 1'b0;  wr_cycle[  575] = 1'b1;  addr_rom[  575]='h00000384;  wr_data_rom[  575]='h000002c5;
    rd_cycle[  576] = 1'b0;  wr_cycle[  576] = 1'b1;  addr_rom[  576]='h00000314;  wr_data_rom[  576]='h000003bb;
    rd_cycle[  577] = 1'b1;  wr_cycle[  577] = 1'b0;  addr_rom[  577]='h00000320;  wr_data_rom[  577]='h00000000;
    rd_cycle[  578] = 1'b1;  wr_cycle[  578] = 1'b0;  addr_rom[  578]='h00000338;  wr_data_rom[  578]='h00000000;
    rd_cycle[  579] = 1'b1;  wr_cycle[  579] = 1'b0;  addr_rom[  579]='h000003ec;  wr_data_rom[  579]='h00000000;
    rd_cycle[  580] = 1'b0;  wr_cycle[  580] = 1'b1;  addr_rom[  580]='h000002a8;  wr_data_rom[  580]='h00000011;
    rd_cycle[  581] = 1'b1;  wr_cycle[  581] = 1'b0;  addr_rom[  581]='h000000e4;  wr_data_rom[  581]='h00000000;
    rd_cycle[  582] = 1'b1;  wr_cycle[  582] = 1'b0;  addr_rom[  582]='h0000003c;  wr_data_rom[  582]='h00000000;
    rd_cycle[  583] = 1'b1;  wr_cycle[  583] = 1'b0;  addr_rom[  583]='h000002ec;  wr_data_rom[  583]='h00000000;
    rd_cycle[  584] = 1'b0;  wr_cycle[  584] = 1'b1;  addr_rom[  584]='h00000380;  wr_data_rom[  584]='h0000022e;
    rd_cycle[  585] = 1'b0;  wr_cycle[  585] = 1'b1;  addr_rom[  585]='h00000178;  wr_data_rom[  585]='h00000134;
    rd_cycle[  586] = 1'b0;  wr_cycle[  586] = 1'b1;  addr_rom[  586]='h0000015c;  wr_data_rom[  586]='h000003f8;
    rd_cycle[  587] = 1'b0;  wr_cycle[  587] = 1'b1;  addr_rom[  587]='h0000005c;  wr_data_rom[  587]='h0000033e;
    rd_cycle[  588] = 1'b0;  wr_cycle[  588] = 1'b1;  addr_rom[  588]='h000001d4;  wr_data_rom[  588]='h00000028;
    rd_cycle[  589] = 1'b0;  wr_cycle[  589] = 1'b1;  addr_rom[  589]='h00000098;  wr_data_rom[  589]='h00000014;
    rd_cycle[  590] = 1'b1;  wr_cycle[  590] = 1'b0;  addr_rom[  590]='h000000c4;  wr_data_rom[  590]='h00000000;
    rd_cycle[  591] = 1'b0;  wr_cycle[  591] = 1'b1;  addr_rom[  591]='h0000016c;  wr_data_rom[  591]='h000000ad;
    rd_cycle[  592] = 1'b1;  wr_cycle[  592] = 1'b0;  addr_rom[  592]='h0000027c;  wr_data_rom[  592]='h00000000;
    rd_cycle[  593] = 1'b0;  wr_cycle[  593] = 1'b1;  addr_rom[  593]='h00000300;  wr_data_rom[  593]='h000000e2;
    rd_cycle[  594] = 1'b1;  wr_cycle[  594] = 1'b0;  addr_rom[  594]='h00000264;  wr_data_rom[  594]='h00000000;
    rd_cycle[  595] = 1'b1;  wr_cycle[  595] = 1'b0;  addr_rom[  595]='h0000017c;  wr_data_rom[  595]='h00000000;
    rd_cycle[  596] = 1'b0;  wr_cycle[  596] = 1'b1;  addr_rom[  596]='h000000e8;  wr_data_rom[  596]='h000000b9;
    rd_cycle[  597] = 1'b0;  wr_cycle[  597] = 1'b1;  addr_rom[  597]='h000002a0;  wr_data_rom[  597]='h00000137;
    rd_cycle[  598] = 1'b1;  wr_cycle[  598] = 1'b0;  addr_rom[  598]='h00000104;  wr_data_rom[  598]='h00000000;
    rd_cycle[  599] = 1'b0;  wr_cycle[  599] = 1'b1;  addr_rom[  599]='h00000118;  wr_data_rom[  599]='h000002ea;
    rd_cycle[  600] = 1'b1;  wr_cycle[  600] = 1'b0;  addr_rom[  600]='h000001a8;  wr_data_rom[  600]='h00000000;
    rd_cycle[  601] = 1'b1;  wr_cycle[  601] = 1'b0;  addr_rom[  601]='h000003e8;  wr_data_rom[  601]='h00000000;
    rd_cycle[  602] = 1'b1;  wr_cycle[  602] = 1'b0;  addr_rom[  602]='h000000e4;  wr_data_rom[  602]='h00000000;
    rd_cycle[  603] = 1'b1;  wr_cycle[  603] = 1'b0;  addr_rom[  603]='h000001b0;  wr_data_rom[  603]='h00000000;
    rd_cycle[  604] = 1'b1;  wr_cycle[  604] = 1'b0;  addr_rom[  604]='h00000278;  wr_data_rom[  604]='h00000000;
    rd_cycle[  605] = 1'b1;  wr_cycle[  605] = 1'b0;  addr_rom[  605]='h00000348;  wr_data_rom[  605]='h00000000;
    rd_cycle[  606] = 1'b0;  wr_cycle[  606] = 1'b1;  addr_rom[  606]='h00000024;  wr_data_rom[  606]='h0000028b;
    rd_cycle[  607] = 1'b1;  wr_cycle[  607] = 1'b0;  addr_rom[  607]='h00000034;  wr_data_rom[  607]='h00000000;
    rd_cycle[  608] = 1'b1;  wr_cycle[  608] = 1'b0;  addr_rom[  608]='h00000330;  wr_data_rom[  608]='h00000000;
    rd_cycle[  609] = 1'b0;  wr_cycle[  609] = 1'b1;  addr_rom[  609]='h000001e4;  wr_data_rom[  609]='h000000d0;
    rd_cycle[  610] = 1'b0;  wr_cycle[  610] = 1'b1;  addr_rom[  610]='h000001a0;  wr_data_rom[  610]='h00000218;
    rd_cycle[  611] = 1'b0;  wr_cycle[  611] = 1'b1;  addr_rom[  611]='h00000298;  wr_data_rom[  611]='h000001a3;
    rd_cycle[  612] = 1'b0;  wr_cycle[  612] = 1'b1;  addr_rom[  612]='h00000064;  wr_data_rom[  612]='h00000042;
    rd_cycle[  613] = 1'b1;  wr_cycle[  613] = 1'b0;  addr_rom[  613]='h00000340;  wr_data_rom[  613]='h00000000;
    rd_cycle[  614] = 1'b0;  wr_cycle[  614] = 1'b1;  addr_rom[  614]='h0000037c;  wr_data_rom[  614]='h000002fa;
    rd_cycle[  615] = 1'b0;  wr_cycle[  615] = 1'b1;  addr_rom[  615]='h0000003c;  wr_data_rom[  615]='h0000001a;
    rd_cycle[  616] = 1'b1;  wr_cycle[  616] = 1'b0;  addr_rom[  616]='h000000f4;  wr_data_rom[  616]='h00000000;
    rd_cycle[  617] = 1'b0;  wr_cycle[  617] = 1'b1;  addr_rom[  617]='h000000cc;  wr_data_rom[  617]='h00000144;
    rd_cycle[  618] = 1'b1;  wr_cycle[  618] = 1'b0;  addr_rom[  618]='h0000024c;  wr_data_rom[  618]='h00000000;
    rd_cycle[  619] = 1'b1;  wr_cycle[  619] = 1'b0;  addr_rom[  619]='h00000210;  wr_data_rom[  619]='h00000000;
    rd_cycle[  620] = 1'b1;  wr_cycle[  620] = 1'b0;  addr_rom[  620]='h0000026c;  wr_data_rom[  620]='h00000000;
    rd_cycle[  621] = 1'b0;  wr_cycle[  621] = 1'b1;  addr_rom[  621]='h000001a0;  wr_data_rom[  621]='h000000b5;
    rd_cycle[  622] = 1'b0;  wr_cycle[  622] = 1'b1;  addr_rom[  622]='h00000060;  wr_data_rom[  622]='h00000388;
    rd_cycle[  623] = 1'b1;  wr_cycle[  623] = 1'b0;  addr_rom[  623]='h00000250;  wr_data_rom[  623]='h00000000;
    rd_cycle[  624] = 1'b0;  wr_cycle[  624] = 1'b1;  addr_rom[  624]='h000002cc;  wr_data_rom[  624]='h000002e7;
    rd_cycle[  625] = 1'b1;  wr_cycle[  625] = 1'b0;  addr_rom[  625]='h00000274;  wr_data_rom[  625]='h00000000;
    rd_cycle[  626] = 1'b1;  wr_cycle[  626] = 1'b0;  addr_rom[  626]='h000000ec;  wr_data_rom[  626]='h00000000;
    rd_cycle[  627] = 1'b0;  wr_cycle[  627] = 1'b1;  addr_rom[  627]='h000000f4;  wr_data_rom[  627]='h00000336;
    rd_cycle[  628] = 1'b0;  wr_cycle[  628] = 1'b1;  addr_rom[  628]='h00000308;  wr_data_rom[  628]='h000001b5;
    rd_cycle[  629] = 1'b1;  wr_cycle[  629] = 1'b0;  addr_rom[  629]='h0000011c;  wr_data_rom[  629]='h00000000;
    rd_cycle[  630] = 1'b1;  wr_cycle[  630] = 1'b0;  addr_rom[  630]='h00000314;  wr_data_rom[  630]='h00000000;
    rd_cycle[  631] = 1'b0;  wr_cycle[  631] = 1'b1;  addr_rom[  631]='h00000094;  wr_data_rom[  631]='h000002b9;
    rd_cycle[  632] = 1'b0;  wr_cycle[  632] = 1'b1;  addr_rom[  632]='h00000020;  wr_data_rom[  632]='h0000033c;
    rd_cycle[  633] = 1'b0;  wr_cycle[  633] = 1'b1;  addr_rom[  633]='h0000018c;  wr_data_rom[  633]='h00000139;
    rd_cycle[  634] = 1'b1;  wr_cycle[  634] = 1'b0;  addr_rom[  634]='h00000000;  wr_data_rom[  634]='h00000000;
    rd_cycle[  635] = 1'b0;  wr_cycle[  635] = 1'b1;  addr_rom[  635]='h00000180;  wr_data_rom[  635]='h000003c2;
    rd_cycle[  636] = 1'b0;  wr_cycle[  636] = 1'b1;  addr_rom[  636]='h0000029c;  wr_data_rom[  636]='h00000140;
    rd_cycle[  637] = 1'b0;  wr_cycle[  637] = 1'b1;  addr_rom[  637]='h0000018c;  wr_data_rom[  637]='h00000031;
    rd_cycle[  638] = 1'b0;  wr_cycle[  638] = 1'b1;  addr_rom[  638]='h000002b8;  wr_data_rom[  638]='h0000012e;
    rd_cycle[  639] = 1'b1;  wr_cycle[  639] = 1'b0;  addr_rom[  639]='h00000330;  wr_data_rom[  639]='h00000000;
    rd_cycle[  640] = 1'b1;  wr_cycle[  640] = 1'b0;  addr_rom[  640]='h000000fc;  wr_data_rom[  640]='h00000000;
    rd_cycle[  641] = 1'b0;  wr_cycle[  641] = 1'b1;  addr_rom[  641]='h00000388;  wr_data_rom[  641]='h00000136;
    rd_cycle[  642] = 1'b0;  wr_cycle[  642] = 1'b1;  addr_rom[  642]='h00000198;  wr_data_rom[  642]='h000001ac;
    rd_cycle[  643] = 1'b1;  wr_cycle[  643] = 1'b0;  addr_rom[  643]='h000003a0;  wr_data_rom[  643]='h00000000;
    rd_cycle[  644] = 1'b1;  wr_cycle[  644] = 1'b0;  addr_rom[  644]='h00000374;  wr_data_rom[  644]='h00000000;
    rd_cycle[  645] = 1'b1;  wr_cycle[  645] = 1'b0;  addr_rom[  645]='h00000224;  wr_data_rom[  645]='h00000000;
    rd_cycle[  646] = 1'b0;  wr_cycle[  646] = 1'b1;  addr_rom[  646]='h00000188;  wr_data_rom[  646]='h0000005c;
    rd_cycle[  647] = 1'b1;  wr_cycle[  647] = 1'b0;  addr_rom[  647]='h000002b0;  wr_data_rom[  647]='h00000000;
    rd_cycle[  648] = 1'b0;  wr_cycle[  648] = 1'b1;  addr_rom[  648]='h00000334;  wr_data_rom[  648]='h000002e2;
    rd_cycle[  649] = 1'b1;  wr_cycle[  649] = 1'b0;  addr_rom[  649]='h000001cc;  wr_data_rom[  649]='h00000000;
    rd_cycle[  650] = 1'b0;  wr_cycle[  650] = 1'b1;  addr_rom[  650]='h0000018c;  wr_data_rom[  650]='h0000034b;
    rd_cycle[  651] = 1'b1;  wr_cycle[  651] = 1'b0;  addr_rom[  651]='h000002e0;  wr_data_rom[  651]='h00000000;
    rd_cycle[  652] = 1'b0;  wr_cycle[  652] = 1'b1;  addr_rom[  652]='h0000022c;  wr_data_rom[  652]='h00000081;
    rd_cycle[  653] = 1'b1;  wr_cycle[  653] = 1'b0;  addr_rom[  653]='h00000030;  wr_data_rom[  653]='h00000000;
    rd_cycle[  654] = 1'b0;  wr_cycle[  654] = 1'b1;  addr_rom[  654]='h00000140;  wr_data_rom[  654]='h000000bd;
    rd_cycle[  655] = 1'b1;  wr_cycle[  655] = 1'b0;  addr_rom[  655]='h00000210;  wr_data_rom[  655]='h00000000;
    rd_cycle[  656] = 1'b1;  wr_cycle[  656] = 1'b0;  addr_rom[  656]='h000000bc;  wr_data_rom[  656]='h00000000;
    rd_cycle[  657] = 1'b0;  wr_cycle[  657] = 1'b1;  addr_rom[  657]='h0000003c;  wr_data_rom[  657]='h000003cc;
    rd_cycle[  658] = 1'b0;  wr_cycle[  658] = 1'b1;  addr_rom[  658]='h000000e4;  wr_data_rom[  658]='h000000bb;
    rd_cycle[  659] = 1'b0;  wr_cycle[  659] = 1'b1;  addr_rom[  659]='h0000032c;  wr_data_rom[  659]='h00000163;
    rd_cycle[  660] = 1'b0;  wr_cycle[  660] = 1'b1;  addr_rom[  660]='h00000280;  wr_data_rom[  660]='h000002bb;
    rd_cycle[  661] = 1'b0;  wr_cycle[  661] = 1'b1;  addr_rom[  661]='h00000118;  wr_data_rom[  661]='h000003e0;
    rd_cycle[  662] = 1'b1;  wr_cycle[  662] = 1'b0;  addr_rom[  662]='h00000044;  wr_data_rom[  662]='h00000000;
    rd_cycle[  663] = 1'b1;  wr_cycle[  663] = 1'b0;  addr_rom[  663]='h0000026c;  wr_data_rom[  663]='h00000000;
    rd_cycle[  664] = 1'b0;  wr_cycle[  664] = 1'b1;  addr_rom[  664]='h00000294;  wr_data_rom[  664]='h00000354;
    rd_cycle[  665] = 1'b1;  wr_cycle[  665] = 1'b0;  addr_rom[  665]='h000000d8;  wr_data_rom[  665]='h00000000;
    rd_cycle[  666] = 1'b0;  wr_cycle[  666] = 1'b1;  addr_rom[  666]='h000003e8;  wr_data_rom[  666]='h00000169;
    rd_cycle[  667] = 1'b1;  wr_cycle[  667] = 1'b0;  addr_rom[  667]='h00000214;  wr_data_rom[  667]='h00000000;
    rd_cycle[  668] = 1'b1;  wr_cycle[  668] = 1'b0;  addr_rom[  668]='h000003c0;  wr_data_rom[  668]='h00000000;
    rd_cycle[  669] = 1'b1;  wr_cycle[  669] = 1'b0;  addr_rom[  669]='h000001dc;  wr_data_rom[  669]='h00000000;
    rd_cycle[  670] = 1'b0;  wr_cycle[  670] = 1'b1;  addr_rom[  670]='h00000398;  wr_data_rom[  670]='h000002fe;
    rd_cycle[  671] = 1'b0;  wr_cycle[  671] = 1'b1;  addr_rom[  671]='h00000244;  wr_data_rom[  671]='h00000159;
    rd_cycle[  672] = 1'b0;  wr_cycle[  672] = 1'b1;  addr_rom[  672]='h00000164;  wr_data_rom[  672]='h000003b7;
    rd_cycle[  673] = 1'b0;  wr_cycle[  673] = 1'b1;  addr_rom[  673]='h000001e0;  wr_data_rom[  673]='h00000105;
    rd_cycle[  674] = 1'b1;  wr_cycle[  674] = 1'b0;  addr_rom[  674]='h00000294;  wr_data_rom[  674]='h00000000;
    rd_cycle[  675] = 1'b1;  wr_cycle[  675] = 1'b0;  addr_rom[  675]='h00000250;  wr_data_rom[  675]='h00000000;
    rd_cycle[  676] = 1'b0;  wr_cycle[  676] = 1'b1;  addr_rom[  676]='h00000308;  wr_data_rom[  676]='h000000f5;
    rd_cycle[  677] = 1'b0;  wr_cycle[  677] = 1'b1;  addr_rom[  677]='h0000014c;  wr_data_rom[  677]='h00000130;
    rd_cycle[  678] = 1'b0;  wr_cycle[  678] = 1'b1;  addr_rom[  678]='h00000390;  wr_data_rom[  678]='h0000023b;
    rd_cycle[  679] = 1'b1;  wr_cycle[  679] = 1'b0;  addr_rom[  679]='h00000148;  wr_data_rom[  679]='h00000000;
    rd_cycle[  680] = 1'b1;  wr_cycle[  680] = 1'b0;  addr_rom[  680]='h000001d0;  wr_data_rom[  680]='h00000000;
    rd_cycle[  681] = 1'b0;  wr_cycle[  681] = 1'b1;  addr_rom[  681]='h000001fc;  wr_data_rom[  681]='h00000182;
    rd_cycle[  682] = 1'b0;  wr_cycle[  682] = 1'b1;  addr_rom[  682]='h00000114;  wr_data_rom[  682]='h000002d0;
    rd_cycle[  683] = 1'b1;  wr_cycle[  683] = 1'b0;  addr_rom[  683]='h00000258;  wr_data_rom[  683]='h00000000;
    rd_cycle[  684] = 1'b1;  wr_cycle[  684] = 1'b0;  addr_rom[  684]='h000001d8;  wr_data_rom[  684]='h00000000;
    rd_cycle[  685] = 1'b0;  wr_cycle[  685] = 1'b1;  addr_rom[  685]='h000003b0;  wr_data_rom[  685]='h00000278;
    rd_cycle[  686] = 1'b0;  wr_cycle[  686] = 1'b1;  addr_rom[  686]='h0000024c;  wr_data_rom[  686]='h000001c5;
    rd_cycle[  687] = 1'b1;  wr_cycle[  687] = 1'b0;  addr_rom[  687]='h000002a4;  wr_data_rom[  687]='h00000000;
    rd_cycle[  688] = 1'b1;  wr_cycle[  688] = 1'b0;  addr_rom[  688]='h000001f8;  wr_data_rom[  688]='h00000000;
    rd_cycle[  689] = 1'b1;  wr_cycle[  689] = 1'b0;  addr_rom[  689]='h000001b4;  wr_data_rom[  689]='h00000000;
    rd_cycle[  690] = 1'b1;  wr_cycle[  690] = 1'b0;  addr_rom[  690]='h000002bc;  wr_data_rom[  690]='h00000000;
    rd_cycle[  691] = 1'b1;  wr_cycle[  691] = 1'b0;  addr_rom[  691]='h00000238;  wr_data_rom[  691]='h00000000;
    rd_cycle[  692] = 1'b1;  wr_cycle[  692] = 1'b0;  addr_rom[  692]='h000003c8;  wr_data_rom[  692]='h00000000;
    rd_cycle[  693] = 1'b0;  wr_cycle[  693] = 1'b1;  addr_rom[  693]='h00000198;  wr_data_rom[  693]='h000001f8;
    rd_cycle[  694] = 1'b1;  wr_cycle[  694] = 1'b0;  addr_rom[  694]='h000001a0;  wr_data_rom[  694]='h00000000;
    rd_cycle[  695] = 1'b1;  wr_cycle[  695] = 1'b0;  addr_rom[  695]='h000002bc;  wr_data_rom[  695]='h00000000;
    rd_cycle[  696] = 1'b1;  wr_cycle[  696] = 1'b0;  addr_rom[  696]='h00000340;  wr_data_rom[  696]='h00000000;
    rd_cycle[  697] = 1'b1;  wr_cycle[  697] = 1'b0;  addr_rom[  697]='h000000b4;  wr_data_rom[  697]='h00000000;
    rd_cycle[  698] = 1'b0;  wr_cycle[  698] = 1'b1;  addr_rom[  698]='h00000348;  wr_data_rom[  698]='h000001c1;
    rd_cycle[  699] = 1'b0;  wr_cycle[  699] = 1'b1;  addr_rom[  699]='h000000a4;  wr_data_rom[  699]='h000002c2;
    rd_cycle[  700] = 1'b1;  wr_cycle[  700] = 1'b0;  addr_rom[  700]='h00000368;  wr_data_rom[  700]='h00000000;
    rd_cycle[  701] = 1'b1;  wr_cycle[  701] = 1'b0;  addr_rom[  701]='h0000009c;  wr_data_rom[  701]='h00000000;
    rd_cycle[  702] = 1'b0;  wr_cycle[  702] = 1'b1;  addr_rom[  702]='h000003d4;  wr_data_rom[  702]='h0000033e;
    rd_cycle[  703] = 1'b0;  wr_cycle[  703] = 1'b1;  addr_rom[  703]='h000002d4;  wr_data_rom[  703]='h0000033c;
    rd_cycle[  704] = 1'b0;  wr_cycle[  704] = 1'b1;  addr_rom[  704]='h00000378;  wr_data_rom[  704]='h00000344;
    rd_cycle[  705] = 1'b1;  wr_cycle[  705] = 1'b0;  addr_rom[  705]='h00000340;  wr_data_rom[  705]='h00000000;
    rd_cycle[  706] = 1'b0;  wr_cycle[  706] = 1'b1;  addr_rom[  706]='h000000cc;  wr_data_rom[  706]='h000000b8;
    rd_cycle[  707] = 1'b1;  wr_cycle[  707] = 1'b0;  addr_rom[  707]='h00000098;  wr_data_rom[  707]='h00000000;
    rd_cycle[  708] = 1'b0;  wr_cycle[  708] = 1'b1;  addr_rom[  708]='h00000074;  wr_data_rom[  708]='h000001b9;
    rd_cycle[  709] = 1'b0;  wr_cycle[  709] = 1'b1;  addr_rom[  709]='h00000228;  wr_data_rom[  709]='h00000062;
    rd_cycle[  710] = 1'b1;  wr_cycle[  710] = 1'b0;  addr_rom[  710]='h00000340;  wr_data_rom[  710]='h00000000;
    rd_cycle[  711] = 1'b0;  wr_cycle[  711] = 1'b1;  addr_rom[  711]='h00000298;  wr_data_rom[  711]='h000000e4;
    rd_cycle[  712] = 1'b1;  wr_cycle[  712] = 1'b0;  addr_rom[  712]='h000002d8;  wr_data_rom[  712]='h00000000;
    rd_cycle[  713] = 1'b1;  wr_cycle[  713] = 1'b0;  addr_rom[  713]='h0000005c;  wr_data_rom[  713]='h00000000;
    rd_cycle[  714] = 1'b0;  wr_cycle[  714] = 1'b1;  addr_rom[  714]='h00000384;  wr_data_rom[  714]='h000000d3;
    rd_cycle[  715] = 1'b0;  wr_cycle[  715] = 1'b1;  addr_rom[  715]='h000003a4;  wr_data_rom[  715]='h0000025f;
    rd_cycle[  716] = 1'b0;  wr_cycle[  716] = 1'b1;  addr_rom[  716]='h000003b0;  wr_data_rom[  716]='h000003ea;
    rd_cycle[  717] = 1'b0;  wr_cycle[  717] = 1'b1;  addr_rom[  717]='h00000040;  wr_data_rom[  717]='h000001d2;
    rd_cycle[  718] = 1'b1;  wr_cycle[  718] = 1'b0;  addr_rom[  718]='h00000130;  wr_data_rom[  718]='h00000000;
    rd_cycle[  719] = 1'b1;  wr_cycle[  719] = 1'b0;  addr_rom[  719]='h000002f4;  wr_data_rom[  719]='h00000000;
    rd_cycle[  720] = 1'b0;  wr_cycle[  720] = 1'b1;  addr_rom[  720]='h000002e4;  wr_data_rom[  720]='h00000168;
    rd_cycle[  721] = 1'b1;  wr_cycle[  721] = 1'b0;  addr_rom[  721]='h000003f4;  wr_data_rom[  721]='h00000000;
    rd_cycle[  722] = 1'b0;  wr_cycle[  722] = 1'b1;  addr_rom[  722]='h00000280;  wr_data_rom[  722]='h000000e0;
    rd_cycle[  723] = 1'b1;  wr_cycle[  723] = 1'b0;  addr_rom[  723]='h0000015c;  wr_data_rom[  723]='h00000000;
    rd_cycle[  724] = 1'b0;  wr_cycle[  724] = 1'b1;  addr_rom[  724]='h000000d0;  wr_data_rom[  724]='h000000a1;
    rd_cycle[  725] = 1'b0;  wr_cycle[  725] = 1'b1;  addr_rom[  725]='h00000168;  wr_data_rom[  725]='h000002c8;
    rd_cycle[  726] = 1'b0;  wr_cycle[  726] = 1'b1;  addr_rom[  726]='h00000318;  wr_data_rom[  726]='h000003a3;
    rd_cycle[  727] = 1'b0;  wr_cycle[  727] = 1'b1;  addr_rom[  727]='h00000050;  wr_data_rom[  727]='h00000041;
    rd_cycle[  728] = 1'b1;  wr_cycle[  728] = 1'b0;  addr_rom[  728]='h000001fc;  wr_data_rom[  728]='h00000000;
    rd_cycle[  729] = 1'b1;  wr_cycle[  729] = 1'b0;  addr_rom[  729]='h000003d0;  wr_data_rom[  729]='h00000000;
    rd_cycle[  730] = 1'b1;  wr_cycle[  730] = 1'b0;  addr_rom[  730]='h0000036c;  wr_data_rom[  730]='h00000000;
    rd_cycle[  731] = 1'b0;  wr_cycle[  731] = 1'b1;  addr_rom[  731]='h0000003c;  wr_data_rom[  731]='h00000332;
    rd_cycle[  732] = 1'b1;  wr_cycle[  732] = 1'b0;  addr_rom[  732]='h00000364;  wr_data_rom[  732]='h00000000;
    rd_cycle[  733] = 1'b1;  wr_cycle[  733] = 1'b0;  addr_rom[  733]='h00000198;  wr_data_rom[  733]='h00000000;
    rd_cycle[  734] = 1'b0;  wr_cycle[  734] = 1'b1;  addr_rom[  734]='h0000028c;  wr_data_rom[  734]='h000003af;
    rd_cycle[  735] = 1'b0;  wr_cycle[  735] = 1'b1;  addr_rom[  735]='h00000164;  wr_data_rom[  735]='h00000159;
    rd_cycle[  736] = 1'b0;  wr_cycle[  736] = 1'b1;  addr_rom[  736]='h000002c8;  wr_data_rom[  736]='h000003d1;
    rd_cycle[  737] = 1'b1;  wr_cycle[  737] = 1'b0;  addr_rom[  737]='h0000017c;  wr_data_rom[  737]='h00000000;
    rd_cycle[  738] = 1'b1;  wr_cycle[  738] = 1'b0;  addr_rom[  738]='h00000008;  wr_data_rom[  738]='h00000000;
    rd_cycle[  739] = 1'b0;  wr_cycle[  739] = 1'b1;  addr_rom[  739]='h000001c0;  wr_data_rom[  739]='h0000036c;
    rd_cycle[  740] = 1'b0;  wr_cycle[  740] = 1'b1;  addr_rom[  740]='h00000100;  wr_data_rom[  740]='h00000079;
    rd_cycle[  741] = 1'b1;  wr_cycle[  741] = 1'b0;  addr_rom[  741]='h00000180;  wr_data_rom[  741]='h00000000;
    rd_cycle[  742] = 1'b1;  wr_cycle[  742] = 1'b0;  addr_rom[  742]='h00000060;  wr_data_rom[  742]='h00000000;
    rd_cycle[  743] = 1'b0;  wr_cycle[  743] = 1'b1;  addr_rom[  743]='h00000228;  wr_data_rom[  743]='h000002a6;
    rd_cycle[  744] = 1'b0;  wr_cycle[  744] = 1'b1;  addr_rom[  744]='h000000c8;  wr_data_rom[  744]='h0000001c;
    rd_cycle[  745] = 1'b1;  wr_cycle[  745] = 1'b0;  addr_rom[  745]='h00000390;  wr_data_rom[  745]='h00000000;
    rd_cycle[  746] = 1'b0;  wr_cycle[  746] = 1'b1;  addr_rom[  746]='h000000ec;  wr_data_rom[  746]='h00000293;
    rd_cycle[  747] = 1'b1;  wr_cycle[  747] = 1'b0;  addr_rom[  747]='h000000f8;  wr_data_rom[  747]='h00000000;
    rd_cycle[  748] = 1'b0;  wr_cycle[  748] = 1'b1;  addr_rom[  748]='h00000004;  wr_data_rom[  748]='h000003c0;
    rd_cycle[  749] = 1'b1;  wr_cycle[  749] = 1'b0;  addr_rom[  749]='h000001bc;  wr_data_rom[  749]='h00000000;
    rd_cycle[  750] = 1'b0;  wr_cycle[  750] = 1'b1;  addr_rom[  750]='h000002c8;  wr_data_rom[  750]='h00000018;
    rd_cycle[  751] = 1'b1;  wr_cycle[  751] = 1'b0;  addr_rom[  751]='h00000348;  wr_data_rom[  751]='h00000000;
    rd_cycle[  752] = 1'b0;  wr_cycle[  752] = 1'b1;  addr_rom[  752]='h00000228;  wr_data_rom[  752]='h00000177;
    rd_cycle[  753] = 1'b0;  wr_cycle[  753] = 1'b1;  addr_rom[  753]='h00000130;  wr_data_rom[  753]='h00000025;
    rd_cycle[  754] = 1'b1;  wr_cycle[  754] = 1'b0;  addr_rom[  754]='h000002d4;  wr_data_rom[  754]='h00000000;
    rd_cycle[  755] = 1'b0;  wr_cycle[  755] = 1'b1;  addr_rom[  755]='h00000394;  wr_data_rom[  755]='h000003db;
    rd_cycle[  756] = 1'b0;  wr_cycle[  756] = 1'b1;  addr_rom[  756]='h0000022c;  wr_data_rom[  756]='h00000141;
    rd_cycle[  757] = 1'b0;  wr_cycle[  757] = 1'b1;  addr_rom[  757]='h00000364;  wr_data_rom[  757]='h0000005c;
    rd_cycle[  758] = 1'b0;  wr_cycle[  758] = 1'b1;  addr_rom[  758]='h0000016c;  wr_data_rom[  758]='h00000385;
    rd_cycle[  759] = 1'b0;  wr_cycle[  759] = 1'b1;  addr_rom[  759]='h000002b8;  wr_data_rom[  759]='h0000030b;
    rd_cycle[  760] = 1'b1;  wr_cycle[  760] = 1'b0;  addr_rom[  760]='h000003c8;  wr_data_rom[  760]='h00000000;
    rd_cycle[  761] = 1'b1;  wr_cycle[  761] = 1'b0;  addr_rom[  761]='h000001f8;  wr_data_rom[  761]='h00000000;
    rd_cycle[  762] = 1'b1;  wr_cycle[  762] = 1'b0;  addr_rom[  762]='h00000014;  wr_data_rom[  762]='h00000000;
    rd_cycle[  763] = 1'b1;  wr_cycle[  763] = 1'b0;  addr_rom[  763]='h0000001c;  wr_data_rom[  763]='h00000000;
    rd_cycle[  764] = 1'b0;  wr_cycle[  764] = 1'b1;  addr_rom[  764]='h000002c4;  wr_data_rom[  764]='h000001dc;
    rd_cycle[  765] = 1'b0;  wr_cycle[  765] = 1'b1;  addr_rom[  765]='h000001d0;  wr_data_rom[  765]='h00000117;
    rd_cycle[  766] = 1'b0;  wr_cycle[  766] = 1'b1;  addr_rom[  766]='h00000160;  wr_data_rom[  766]='h0000033a;
    rd_cycle[  767] = 1'b0;  wr_cycle[  767] = 1'b1;  addr_rom[  767]='h00000288;  wr_data_rom[  767]='h000003ef;
    rd_cycle[  768] = 1'b0;  wr_cycle[  768] = 1'b1;  addr_rom[  768]='h0000031c;  wr_data_rom[  768]='h00000391;
    rd_cycle[  769] = 1'b0;  wr_cycle[  769] = 1'b1;  addr_rom[  769]='h00000024;  wr_data_rom[  769]='h0000005f;
    rd_cycle[  770] = 1'b1;  wr_cycle[  770] = 1'b0;  addr_rom[  770]='h0000008c;  wr_data_rom[  770]='h00000000;
    rd_cycle[  771] = 1'b1;  wr_cycle[  771] = 1'b0;  addr_rom[  771]='h00000224;  wr_data_rom[  771]='h00000000;
    rd_cycle[  772] = 1'b1;  wr_cycle[  772] = 1'b0;  addr_rom[  772]='h000002b8;  wr_data_rom[  772]='h00000000;
    rd_cycle[  773] = 1'b0;  wr_cycle[  773] = 1'b1;  addr_rom[  773]='h00000168;  wr_data_rom[  773]='h00000082;
    rd_cycle[  774] = 1'b1;  wr_cycle[  774] = 1'b0;  addr_rom[  774]='h00000134;  wr_data_rom[  774]='h00000000;
    rd_cycle[  775] = 1'b0;  wr_cycle[  775] = 1'b1;  addr_rom[  775]='h00000034;  wr_data_rom[  775]='h00000308;
    rd_cycle[  776] = 1'b1;  wr_cycle[  776] = 1'b0;  addr_rom[  776]='h0000029c;  wr_data_rom[  776]='h00000000;
    rd_cycle[  777] = 1'b0;  wr_cycle[  777] = 1'b1;  addr_rom[  777]='h00000154;  wr_data_rom[  777]='h00000233;
    rd_cycle[  778] = 1'b0;  wr_cycle[  778] = 1'b1;  addr_rom[  778]='h00000164;  wr_data_rom[  778]='h000001eb;
    rd_cycle[  779] = 1'b0;  wr_cycle[  779] = 1'b1;  addr_rom[  779]='h00000080;  wr_data_rom[  779]='h00000192;
    rd_cycle[  780] = 1'b0;  wr_cycle[  780] = 1'b1;  addr_rom[  780]='h0000008c;  wr_data_rom[  780]='h00000095;
    rd_cycle[  781] = 1'b1;  wr_cycle[  781] = 1'b0;  addr_rom[  781]='h00000144;  wr_data_rom[  781]='h00000000;
    rd_cycle[  782] = 1'b1;  wr_cycle[  782] = 1'b0;  addr_rom[  782]='h0000022c;  wr_data_rom[  782]='h00000000;
    rd_cycle[  783] = 1'b1;  wr_cycle[  783] = 1'b0;  addr_rom[  783]='h00000290;  wr_data_rom[  783]='h00000000;
    rd_cycle[  784] = 1'b0;  wr_cycle[  784] = 1'b1;  addr_rom[  784]='h000001b8;  wr_data_rom[  784]='h000001eb;
    rd_cycle[  785] = 1'b1;  wr_cycle[  785] = 1'b0;  addr_rom[  785]='h000000dc;  wr_data_rom[  785]='h00000000;
    rd_cycle[  786] = 1'b1;  wr_cycle[  786] = 1'b0;  addr_rom[  786]='h000000e0;  wr_data_rom[  786]='h00000000;
    rd_cycle[  787] = 1'b1;  wr_cycle[  787] = 1'b0;  addr_rom[  787]='h00000050;  wr_data_rom[  787]='h00000000;
    rd_cycle[  788] = 1'b0;  wr_cycle[  788] = 1'b1;  addr_rom[  788]='h00000308;  wr_data_rom[  788]='h0000035d;
    rd_cycle[  789] = 1'b0;  wr_cycle[  789] = 1'b1;  addr_rom[  789]='h00000390;  wr_data_rom[  789]='h000002dc;
    rd_cycle[  790] = 1'b0;  wr_cycle[  790] = 1'b1;  addr_rom[  790]='h0000026c;  wr_data_rom[  790]='h0000038b;
    rd_cycle[  791] = 1'b0;  wr_cycle[  791] = 1'b1;  addr_rom[  791]='h000001f4;  wr_data_rom[  791]='h00000279;
    rd_cycle[  792] = 1'b0;  wr_cycle[  792] = 1'b1;  addr_rom[  792]='h00000264;  wr_data_rom[  792]='h000002f7;
    rd_cycle[  793] = 1'b1;  wr_cycle[  793] = 1'b0;  addr_rom[  793]='h00000078;  wr_data_rom[  793]='h00000000;
    rd_cycle[  794] = 1'b1;  wr_cycle[  794] = 1'b0;  addr_rom[  794]='h000003c8;  wr_data_rom[  794]='h00000000;
    rd_cycle[  795] = 1'b0;  wr_cycle[  795] = 1'b1;  addr_rom[  795]='h00000124;  wr_data_rom[  795]='h000001b8;
    rd_cycle[  796] = 1'b0;  wr_cycle[  796] = 1'b1;  addr_rom[  796]='h000002d4;  wr_data_rom[  796]='h00000238;
    rd_cycle[  797] = 1'b0;  wr_cycle[  797] = 1'b1;  addr_rom[  797]='h00000238;  wr_data_rom[  797]='h00000357;
    rd_cycle[  798] = 1'b1;  wr_cycle[  798] = 1'b0;  addr_rom[  798]='h00000380;  wr_data_rom[  798]='h00000000;
    rd_cycle[  799] = 1'b1;  wr_cycle[  799] = 1'b0;  addr_rom[  799]='h0000007c;  wr_data_rom[  799]='h00000000;
    rd_cycle[  800] = 1'b1;  wr_cycle[  800] = 1'b0;  addr_rom[  800]='h00000154;  wr_data_rom[  800]='h00000000;
    rd_cycle[  801] = 1'b0;  wr_cycle[  801] = 1'b1;  addr_rom[  801]='h000000f0;  wr_data_rom[  801]='h00000261;
    rd_cycle[  802] = 1'b0;  wr_cycle[  802] = 1'b1;  addr_rom[  802]='h000003dc;  wr_data_rom[  802]='h0000036e;
    rd_cycle[  803] = 1'b0;  wr_cycle[  803] = 1'b1;  addr_rom[  803]='h000001e8;  wr_data_rom[  803]='h00000058;
    rd_cycle[  804] = 1'b0;  wr_cycle[  804] = 1'b1;  addr_rom[  804]='h00000090;  wr_data_rom[  804]='h00000220;
    rd_cycle[  805] = 1'b1;  wr_cycle[  805] = 1'b0;  addr_rom[  805]='h000003c8;  wr_data_rom[  805]='h00000000;
    rd_cycle[  806] = 1'b0;  wr_cycle[  806] = 1'b1;  addr_rom[  806]='h000003e0;  wr_data_rom[  806]='h00000093;
    rd_cycle[  807] = 1'b0;  wr_cycle[  807] = 1'b1;  addr_rom[  807]='h00000234;  wr_data_rom[  807]='h000000d9;
    rd_cycle[  808] = 1'b0;  wr_cycle[  808] = 1'b1;  addr_rom[  808]='h000000b8;  wr_data_rom[  808]='h000002f6;
    rd_cycle[  809] = 1'b1;  wr_cycle[  809] = 1'b0;  addr_rom[  809]='h000002f0;  wr_data_rom[  809]='h00000000;
    rd_cycle[  810] = 1'b0;  wr_cycle[  810] = 1'b1;  addr_rom[  810]='h00000088;  wr_data_rom[  810]='h000000ca;
    rd_cycle[  811] = 1'b0;  wr_cycle[  811] = 1'b1;  addr_rom[  811]='h00000258;  wr_data_rom[  811]='h000001a1;
    rd_cycle[  812] = 1'b0;  wr_cycle[  812] = 1'b1;  addr_rom[  812]='h00000030;  wr_data_rom[  812]='h000000ac;
    rd_cycle[  813] = 1'b1;  wr_cycle[  813] = 1'b0;  addr_rom[  813]='h000000e4;  wr_data_rom[  813]='h00000000;
    rd_cycle[  814] = 1'b1;  wr_cycle[  814] = 1'b0;  addr_rom[  814]='h00000138;  wr_data_rom[  814]='h00000000;
    rd_cycle[  815] = 1'b0;  wr_cycle[  815] = 1'b1;  addr_rom[  815]='h00000360;  wr_data_rom[  815]='h00000334;
    rd_cycle[  816] = 1'b1;  wr_cycle[  816] = 1'b0;  addr_rom[  816]='h000002ec;  wr_data_rom[  816]='h00000000;
    rd_cycle[  817] = 1'b1;  wr_cycle[  817] = 1'b0;  addr_rom[  817]='h00000370;  wr_data_rom[  817]='h00000000;
    rd_cycle[  818] = 1'b0;  wr_cycle[  818] = 1'b1;  addr_rom[  818]='h0000032c;  wr_data_rom[  818]='h0000022c;
    rd_cycle[  819] = 1'b1;  wr_cycle[  819] = 1'b0;  addr_rom[  819]='h000000b8;  wr_data_rom[  819]='h00000000;
    rd_cycle[  820] = 1'b1;  wr_cycle[  820] = 1'b0;  addr_rom[  820]='h000000a4;  wr_data_rom[  820]='h00000000;
    rd_cycle[  821] = 1'b1;  wr_cycle[  821] = 1'b0;  addr_rom[  821]='h0000016c;  wr_data_rom[  821]='h00000000;
    rd_cycle[  822] = 1'b0;  wr_cycle[  822] = 1'b1;  addr_rom[  822]='h000000e8;  wr_data_rom[  822]='h0000009b;
    rd_cycle[  823] = 1'b0;  wr_cycle[  823] = 1'b1;  addr_rom[  823]='h000003ec;  wr_data_rom[  823]='h00000153;
    rd_cycle[  824] = 1'b0;  wr_cycle[  824] = 1'b1;  addr_rom[  824]='h000000f4;  wr_data_rom[  824]='h0000036f;
    rd_cycle[  825] = 1'b1;  wr_cycle[  825] = 1'b0;  addr_rom[  825]='h0000025c;  wr_data_rom[  825]='h00000000;
    rd_cycle[  826] = 1'b0;  wr_cycle[  826] = 1'b1;  addr_rom[  826]='h0000021c;  wr_data_rom[  826]='h000003f9;
    rd_cycle[  827] = 1'b0;  wr_cycle[  827] = 1'b1;  addr_rom[  827]='h00000228;  wr_data_rom[  827]='h0000031d;
    rd_cycle[  828] = 1'b1;  wr_cycle[  828] = 1'b0;  addr_rom[  828]='h00000298;  wr_data_rom[  828]='h00000000;
    rd_cycle[  829] = 1'b0;  wr_cycle[  829] = 1'b1;  addr_rom[  829]='h0000038c;  wr_data_rom[  829]='h0000035c;
    rd_cycle[  830] = 1'b1;  wr_cycle[  830] = 1'b0;  addr_rom[  830]='h00000150;  wr_data_rom[  830]='h00000000;
    rd_cycle[  831] = 1'b1;  wr_cycle[  831] = 1'b0;  addr_rom[  831]='h000001f4;  wr_data_rom[  831]='h00000000;
    rd_cycle[  832] = 1'b0;  wr_cycle[  832] = 1'b1;  addr_rom[  832]='h000002cc;  wr_data_rom[  832]='h00000088;
    rd_cycle[  833] = 1'b1;  wr_cycle[  833] = 1'b0;  addr_rom[  833]='h00000114;  wr_data_rom[  833]='h00000000;
    rd_cycle[  834] = 1'b1;  wr_cycle[  834] = 1'b0;  addr_rom[  834]='h000003c0;  wr_data_rom[  834]='h00000000;
    rd_cycle[  835] = 1'b1;  wr_cycle[  835] = 1'b0;  addr_rom[  835]='h000002dc;  wr_data_rom[  835]='h00000000;
    rd_cycle[  836] = 1'b1;  wr_cycle[  836] = 1'b0;  addr_rom[  836]='h00000300;  wr_data_rom[  836]='h00000000;
    rd_cycle[  837] = 1'b1;  wr_cycle[  837] = 1'b0;  addr_rom[  837]='h00000104;  wr_data_rom[  837]='h00000000;
    rd_cycle[  838] = 1'b1;  wr_cycle[  838] = 1'b0;  addr_rom[  838]='h000003e4;  wr_data_rom[  838]='h00000000;
    rd_cycle[  839] = 1'b0;  wr_cycle[  839] = 1'b1;  addr_rom[  839]='h00000048;  wr_data_rom[  839]='h00000231;
    rd_cycle[  840] = 1'b1;  wr_cycle[  840] = 1'b0;  addr_rom[  840]='h00000268;  wr_data_rom[  840]='h00000000;
    rd_cycle[  841] = 1'b1;  wr_cycle[  841] = 1'b0;  addr_rom[  841]='h000003d0;  wr_data_rom[  841]='h00000000;
    rd_cycle[  842] = 1'b0;  wr_cycle[  842] = 1'b1;  addr_rom[  842]='h000002f4;  wr_data_rom[  842]='h0000006e;
    rd_cycle[  843] = 1'b0;  wr_cycle[  843] = 1'b1;  addr_rom[  843]='h000001c0;  wr_data_rom[  843]='h00000379;
    rd_cycle[  844] = 1'b1;  wr_cycle[  844] = 1'b0;  addr_rom[  844]='h00000208;  wr_data_rom[  844]='h00000000;
    rd_cycle[  845] = 1'b1;  wr_cycle[  845] = 1'b0;  addr_rom[  845]='h000002ec;  wr_data_rom[  845]='h00000000;
    rd_cycle[  846] = 1'b1;  wr_cycle[  846] = 1'b0;  addr_rom[  846]='h000002d8;  wr_data_rom[  846]='h00000000;
    rd_cycle[  847] = 1'b0;  wr_cycle[  847] = 1'b1;  addr_rom[  847]='h000002e4;  wr_data_rom[  847]='h000002ac;
    rd_cycle[  848] = 1'b1;  wr_cycle[  848] = 1'b0;  addr_rom[  848]='h000001c8;  wr_data_rom[  848]='h00000000;
    rd_cycle[  849] = 1'b0;  wr_cycle[  849] = 1'b1;  addr_rom[  849]='h00000228;  wr_data_rom[  849]='h0000017d;
    rd_cycle[  850] = 1'b0;  wr_cycle[  850] = 1'b1;  addr_rom[  850]='h00000020;  wr_data_rom[  850]='h00000044;
    rd_cycle[  851] = 1'b0;  wr_cycle[  851] = 1'b1;  addr_rom[  851]='h00000020;  wr_data_rom[  851]='h00000157;
    rd_cycle[  852] = 1'b1;  wr_cycle[  852] = 1'b0;  addr_rom[  852]='h000001c4;  wr_data_rom[  852]='h00000000;
    rd_cycle[  853] = 1'b1;  wr_cycle[  853] = 1'b0;  addr_rom[  853]='h000001f8;  wr_data_rom[  853]='h00000000;
    rd_cycle[  854] = 1'b0;  wr_cycle[  854] = 1'b1;  addr_rom[  854]='h00000320;  wr_data_rom[  854]='h00000395;
    rd_cycle[  855] = 1'b1;  wr_cycle[  855] = 1'b0;  addr_rom[  855]='h00000388;  wr_data_rom[  855]='h00000000;
    rd_cycle[  856] = 1'b0;  wr_cycle[  856] = 1'b1;  addr_rom[  856]='h00000268;  wr_data_rom[  856]='h0000001f;
    rd_cycle[  857] = 1'b0;  wr_cycle[  857] = 1'b1;  addr_rom[  857]='h000003c4;  wr_data_rom[  857]='h00000033;
    rd_cycle[  858] = 1'b0;  wr_cycle[  858] = 1'b1;  addr_rom[  858]='h000001b0;  wr_data_rom[  858]='h000003fd;
    rd_cycle[  859] = 1'b0;  wr_cycle[  859] = 1'b1;  addr_rom[  859]='h00000190;  wr_data_rom[  859]='h00000059;
    rd_cycle[  860] = 1'b1;  wr_cycle[  860] = 1'b0;  addr_rom[  860]='h000003f4;  wr_data_rom[  860]='h00000000;
    rd_cycle[  861] = 1'b0;  wr_cycle[  861] = 1'b1;  addr_rom[  861]='h000003f8;  wr_data_rom[  861]='h000002c0;
    rd_cycle[  862] = 1'b0;  wr_cycle[  862] = 1'b1;  addr_rom[  862]='h000001c8;  wr_data_rom[  862]='h00000366;
    rd_cycle[  863] = 1'b0;  wr_cycle[  863] = 1'b1;  addr_rom[  863]='h000001ec;  wr_data_rom[  863]='h0000034e;
    rd_cycle[  864] = 1'b1;  wr_cycle[  864] = 1'b0;  addr_rom[  864]='h00000158;  wr_data_rom[  864]='h00000000;
    rd_cycle[  865] = 1'b1;  wr_cycle[  865] = 1'b0;  addr_rom[  865]='h000003f4;  wr_data_rom[  865]='h00000000;
    rd_cycle[  866] = 1'b1;  wr_cycle[  866] = 1'b0;  addr_rom[  866]='h000003d4;  wr_data_rom[  866]='h00000000;
    rd_cycle[  867] = 1'b0;  wr_cycle[  867] = 1'b1;  addr_rom[  867]='h00000188;  wr_data_rom[  867]='h00000053;
    rd_cycle[  868] = 1'b0;  wr_cycle[  868] = 1'b1;  addr_rom[  868]='h000003e0;  wr_data_rom[  868]='h000001e3;
    rd_cycle[  869] = 1'b1;  wr_cycle[  869] = 1'b0;  addr_rom[  869]='h000003a0;  wr_data_rom[  869]='h00000000;
    rd_cycle[  870] = 1'b0;  wr_cycle[  870] = 1'b1;  addr_rom[  870]='h00000398;  wr_data_rom[  870]='h0000014f;
    rd_cycle[  871] = 1'b1;  wr_cycle[  871] = 1'b0;  addr_rom[  871]='h00000114;  wr_data_rom[  871]='h00000000;
    rd_cycle[  872] = 1'b0;  wr_cycle[  872] = 1'b1;  addr_rom[  872]='h00000248;  wr_data_rom[  872]='h000000a4;
    rd_cycle[  873] = 1'b0;  wr_cycle[  873] = 1'b1;  addr_rom[  873]='h0000016c;  wr_data_rom[  873]='h000000ea;
    rd_cycle[  874] = 1'b1;  wr_cycle[  874] = 1'b0;  addr_rom[  874]='h000001ac;  wr_data_rom[  874]='h00000000;
    rd_cycle[  875] = 1'b1;  wr_cycle[  875] = 1'b0;  addr_rom[  875]='h0000037c;  wr_data_rom[  875]='h00000000;
    rd_cycle[  876] = 1'b1;  wr_cycle[  876] = 1'b0;  addr_rom[  876]='h00000250;  wr_data_rom[  876]='h00000000;
    rd_cycle[  877] = 1'b1;  wr_cycle[  877] = 1'b0;  addr_rom[  877]='h00000180;  wr_data_rom[  877]='h00000000;
    rd_cycle[  878] = 1'b1;  wr_cycle[  878] = 1'b0;  addr_rom[  878]='h000000d0;  wr_data_rom[  878]='h00000000;
    rd_cycle[  879] = 1'b1;  wr_cycle[  879] = 1'b0;  addr_rom[  879]='h00000294;  wr_data_rom[  879]='h00000000;
    rd_cycle[  880] = 1'b0;  wr_cycle[  880] = 1'b1;  addr_rom[  880]='h00000238;  wr_data_rom[  880]='h000003f0;
    rd_cycle[  881] = 1'b1;  wr_cycle[  881] = 1'b0;  addr_rom[  881]='h00000360;  wr_data_rom[  881]='h00000000;
    rd_cycle[  882] = 1'b1;  wr_cycle[  882] = 1'b0;  addr_rom[  882]='h0000010c;  wr_data_rom[  882]='h00000000;
    rd_cycle[  883] = 1'b0;  wr_cycle[  883] = 1'b1;  addr_rom[  883]='h000001f8;  wr_data_rom[  883]='h0000018b;
    rd_cycle[  884] = 1'b0;  wr_cycle[  884] = 1'b1;  addr_rom[  884]='h000003e8;  wr_data_rom[  884]='h000000a0;
    rd_cycle[  885] = 1'b1;  wr_cycle[  885] = 1'b0;  addr_rom[  885]='h000002dc;  wr_data_rom[  885]='h00000000;
    rd_cycle[  886] = 1'b1;  wr_cycle[  886] = 1'b0;  addr_rom[  886]='h00000214;  wr_data_rom[  886]='h00000000;
    rd_cycle[  887] = 1'b1;  wr_cycle[  887] = 1'b0;  addr_rom[  887]='h000002b8;  wr_data_rom[  887]='h00000000;
    rd_cycle[  888] = 1'b0;  wr_cycle[  888] = 1'b1;  addr_rom[  888]='h00000128;  wr_data_rom[  888]='h00000325;
    rd_cycle[  889] = 1'b0;  wr_cycle[  889] = 1'b1;  addr_rom[  889]='h00000108;  wr_data_rom[  889]='h0000003e;
    rd_cycle[  890] = 1'b1;  wr_cycle[  890] = 1'b0;  addr_rom[  890]='h00000224;  wr_data_rom[  890]='h00000000;
    rd_cycle[  891] = 1'b1;  wr_cycle[  891] = 1'b0;  addr_rom[  891]='h00000368;  wr_data_rom[  891]='h00000000;
    rd_cycle[  892] = 1'b0;  wr_cycle[  892] = 1'b1;  addr_rom[  892]='h00000360;  wr_data_rom[  892]='h00000325;
    rd_cycle[  893] = 1'b1;  wr_cycle[  893] = 1'b0;  addr_rom[  893]='h0000005c;  wr_data_rom[  893]='h00000000;
    rd_cycle[  894] = 1'b0;  wr_cycle[  894] = 1'b1;  addr_rom[  894]='h00000388;  wr_data_rom[  894]='h000003e6;
    rd_cycle[  895] = 1'b1;  wr_cycle[  895] = 1'b0;  addr_rom[  895]='h00000030;  wr_data_rom[  895]='h00000000;
    rd_cycle[  896] = 1'b1;  wr_cycle[  896] = 1'b0;  addr_rom[  896]='h00000130;  wr_data_rom[  896]='h00000000;
    rd_cycle[  897] = 1'b1;  wr_cycle[  897] = 1'b0;  addr_rom[  897]='h000002f4;  wr_data_rom[  897]='h00000000;
    rd_cycle[  898] = 1'b1;  wr_cycle[  898] = 1'b0;  addr_rom[  898]='h000002f4;  wr_data_rom[  898]='h00000000;
    rd_cycle[  899] = 1'b1;  wr_cycle[  899] = 1'b0;  addr_rom[  899]='h00000078;  wr_data_rom[  899]='h00000000;
    rd_cycle[  900] = 1'b1;  wr_cycle[  900] = 1'b0;  addr_rom[  900]='h00000150;  wr_data_rom[  900]='h00000000;
    rd_cycle[  901] = 1'b1;  wr_cycle[  901] = 1'b0;  addr_rom[  901]='h00000368;  wr_data_rom[  901]='h00000000;
    rd_cycle[  902] = 1'b1;  wr_cycle[  902] = 1'b0;  addr_rom[  902]='h000001fc;  wr_data_rom[  902]='h00000000;
    rd_cycle[  903] = 1'b0;  wr_cycle[  903] = 1'b1;  addr_rom[  903]='h0000012c;  wr_data_rom[  903]='h00000163;
    rd_cycle[  904] = 1'b0;  wr_cycle[  904] = 1'b1;  addr_rom[  904]='h00000280;  wr_data_rom[  904]='h00000074;
    rd_cycle[  905] = 1'b0;  wr_cycle[  905] = 1'b1;  addr_rom[  905]='h000002a0;  wr_data_rom[  905]='h000003f4;
    rd_cycle[  906] = 1'b0;  wr_cycle[  906] = 1'b1;  addr_rom[  906]='h000003c4;  wr_data_rom[  906]='h0000007b;
    rd_cycle[  907] = 1'b1;  wr_cycle[  907] = 1'b0;  addr_rom[  907]='h000003bc;  wr_data_rom[  907]='h00000000;
    rd_cycle[  908] = 1'b0;  wr_cycle[  908] = 1'b1;  addr_rom[  908]='h00000158;  wr_data_rom[  908]='h0000036c;
    rd_cycle[  909] = 1'b1;  wr_cycle[  909] = 1'b0;  addr_rom[  909]='h0000010c;  wr_data_rom[  909]='h00000000;
    rd_cycle[  910] = 1'b0;  wr_cycle[  910] = 1'b1;  addr_rom[  910]='h00000168;  wr_data_rom[  910]='h00000052;
    rd_cycle[  911] = 1'b0;  wr_cycle[  911] = 1'b1;  addr_rom[  911]='h000000d0;  wr_data_rom[  911]='h00000240;
    rd_cycle[  912] = 1'b0;  wr_cycle[  912] = 1'b1;  addr_rom[  912]='h000000f8;  wr_data_rom[  912]='h000002c2;
    rd_cycle[  913] = 1'b1;  wr_cycle[  913] = 1'b0;  addr_rom[  913]='h00000110;  wr_data_rom[  913]='h00000000;
    rd_cycle[  914] = 1'b0;  wr_cycle[  914] = 1'b1;  addr_rom[  914]='h00000130;  wr_data_rom[  914]='h0000000e;
    rd_cycle[  915] = 1'b0;  wr_cycle[  915] = 1'b1;  addr_rom[  915]='h00000344;  wr_data_rom[  915]='h00000105;
    rd_cycle[  916] = 1'b1;  wr_cycle[  916] = 1'b0;  addr_rom[  916]='h0000007c;  wr_data_rom[  916]='h00000000;
    rd_cycle[  917] = 1'b0;  wr_cycle[  917] = 1'b1;  addr_rom[  917]='h000000a0;  wr_data_rom[  917]='h0000013c;
    rd_cycle[  918] = 1'b1;  wr_cycle[  918] = 1'b0;  addr_rom[  918]='h00000234;  wr_data_rom[  918]='h00000000;
    rd_cycle[  919] = 1'b1;  wr_cycle[  919] = 1'b0;  addr_rom[  919]='h00000340;  wr_data_rom[  919]='h00000000;
    rd_cycle[  920] = 1'b1;  wr_cycle[  920] = 1'b0;  addr_rom[  920]='h000002cc;  wr_data_rom[  920]='h00000000;
    rd_cycle[  921] = 1'b0;  wr_cycle[  921] = 1'b1;  addr_rom[  921]='h0000038c;  wr_data_rom[  921]='h00000383;
    rd_cycle[  922] = 1'b1;  wr_cycle[  922] = 1'b0;  addr_rom[  922]='h000002d4;  wr_data_rom[  922]='h00000000;
    rd_cycle[  923] = 1'b0;  wr_cycle[  923] = 1'b1;  addr_rom[  923]='h00000274;  wr_data_rom[  923]='h00000071;
    rd_cycle[  924] = 1'b1;  wr_cycle[  924] = 1'b0;  addr_rom[  924]='h00000240;  wr_data_rom[  924]='h00000000;
    rd_cycle[  925] = 1'b1;  wr_cycle[  925] = 1'b0;  addr_rom[  925]='h00000014;  wr_data_rom[  925]='h00000000;
    rd_cycle[  926] = 1'b1;  wr_cycle[  926] = 1'b0;  addr_rom[  926]='h00000290;  wr_data_rom[  926]='h00000000;
    rd_cycle[  927] = 1'b0;  wr_cycle[  927] = 1'b1;  addr_rom[  927]='h00000080;  wr_data_rom[  927]='h000000af;
    rd_cycle[  928] = 1'b0;  wr_cycle[  928] = 1'b1;  addr_rom[  928]='h0000019c;  wr_data_rom[  928]='h000003d5;
    rd_cycle[  929] = 1'b0;  wr_cycle[  929] = 1'b1;  addr_rom[  929]='h000000d0;  wr_data_rom[  929]='h000001f5;
    rd_cycle[  930] = 1'b0;  wr_cycle[  930] = 1'b1;  addr_rom[  930]='h00000218;  wr_data_rom[  930]='h00000266;
    rd_cycle[  931] = 1'b0;  wr_cycle[  931] = 1'b1;  addr_rom[  931]='h000003f4;  wr_data_rom[  931]='h000000ce;
    rd_cycle[  932] = 1'b1;  wr_cycle[  932] = 1'b0;  addr_rom[  932]='h0000008c;  wr_data_rom[  932]='h00000000;
    rd_cycle[  933] = 1'b0;  wr_cycle[  933] = 1'b1;  addr_rom[  933]='h0000000c;  wr_data_rom[  933]='h0000018b;
    rd_cycle[  934] = 1'b0;  wr_cycle[  934] = 1'b1;  addr_rom[  934]='h000003c4;  wr_data_rom[  934]='h00000391;
    rd_cycle[  935] = 1'b1;  wr_cycle[  935] = 1'b0;  addr_rom[  935]='h0000007c;  wr_data_rom[  935]='h00000000;
    rd_cycle[  936] = 1'b1;  wr_cycle[  936] = 1'b0;  addr_rom[  936]='h00000190;  wr_data_rom[  936]='h00000000;
    rd_cycle[  937] = 1'b1;  wr_cycle[  937] = 1'b0;  addr_rom[  937]='h00000220;  wr_data_rom[  937]='h00000000;
    rd_cycle[  938] = 1'b1;  wr_cycle[  938] = 1'b0;  addr_rom[  938]='h00000198;  wr_data_rom[  938]='h00000000;
    rd_cycle[  939] = 1'b1;  wr_cycle[  939] = 1'b0;  addr_rom[  939]='h000003b4;  wr_data_rom[  939]='h00000000;
    rd_cycle[  940] = 1'b1;  wr_cycle[  940] = 1'b0;  addr_rom[  940]='h000003b4;  wr_data_rom[  940]='h00000000;
    rd_cycle[  941] = 1'b0;  wr_cycle[  941] = 1'b1;  addr_rom[  941]='h00000254;  wr_data_rom[  941]='h000001a1;
    rd_cycle[  942] = 1'b1;  wr_cycle[  942] = 1'b0;  addr_rom[  942]='h00000334;  wr_data_rom[  942]='h00000000;
    rd_cycle[  943] = 1'b0;  wr_cycle[  943] = 1'b1;  addr_rom[  943]='h00000104;  wr_data_rom[  943]='h000001a2;
    rd_cycle[  944] = 1'b1;  wr_cycle[  944] = 1'b0;  addr_rom[  944]='h00000004;  wr_data_rom[  944]='h00000000;
    rd_cycle[  945] = 1'b1;  wr_cycle[  945] = 1'b0;  addr_rom[  945]='h00000350;  wr_data_rom[  945]='h00000000;
    rd_cycle[  946] = 1'b1;  wr_cycle[  946] = 1'b0;  addr_rom[  946]='h000003fc;  wr_data_rom[  946]='h00000000;
    rd_cycle[  947] = 1'b1;  wr_cycle[  947] = 1'b0;  addr_rom[  947]='h00000138;  wr_data_rom[  947]='h00000000;
    rd_cycle[  948] = 1'b0;  wr_cycle[  948] = 1'b1;  addr_rom[  948]='h0000010c;  wr_data_rom[  948]='h00000209;
    rd_cycle[  949] = 1'b1;  wr_cycle[  949] = 1'b0;  addr_rom[  949]='h00000214;  wr_data_rom[  949]='h00000000;
    rd_cycle[  950] = 1'b0;  wr_cycle[  950] = 1'b1;  addr_rom[  950]='h00000390;  wr_data_rom[  950]='h000000e1;
    rd_cycle[  951] = 1'b1;  wr_cycle[  951] = 1'b0;  addr_rom[  951]='h00000184;  wr_data_rom[  951]='h00000000;
    rd_cycle[  952] = 1'b1;  wr_cycle[  952] = 1'b0;  addr_rom[  952]='h000003a4;  wr_data_rom[  952]='h00000000;
    rd_cycle[  953] = 1'b1;  wr_cycle[  953] = 1'b0;  addr_rom[  953]='h00000170;  wr_data_rom[  953]='h00000000;
    rd_cycle[  954] = 1'b1;  wr_cycle[  954] = 1'b0;  addr_rom[  954]='h000001d8;  wr_data_rom[  954]='h00000000;
    rd_cycle[  955] = 1'b0;  wr_cycle[  955] = 1'b1;  addr_rom[  955]='h000002b8;  wr_data_rom[  955]='h000002d9;
    rd_cycle[  956] = 1'b0;  wr_cycle[  956] = 1'b1;  addr_rom[  956]='h000003c0;  wr_data_rom[  956]='h0000024f;
    rd_cycle[  957] = 1'b0;  wr_cycle[  957] = 1'b1;  addr_rom[  957]='h00000018;  wr_data_rom[  957]='h00000262;
    rd_cycle[  958] = 1'b1;  wr_cycle[  958] = 1'b0;  addr_rom[  958]='h000000d0;  wr_data_rom[  958]='h00000000;
    rd_cycle[  959] = 1'b1;  wr_cycle[  959] = 1'b0;  addr_rom[  959]='h00000054;  wr_data_rom[  959]='h00000000;
    rd_cycle[  960] = 1'b1;  wr_cycle[  960] = 1'b0;  addr_rom[  960]='h000000e0;  wr_data_rom[  960]='h00000000;
    rd_cycle[  961] = 1'b0;  wr_cycle[  961] = 1'b1;  addr_rom[  961]='h000003f8;  wr_data_rom[  961]='h00000291;
    rd_cycle[  962] = 1'b1;  wr_cycle[  962] = 1'b0;  addr_rom[  962]='h00000160;  wr_data_rom[  962]='h00000000;
    rd_cycle[  963] = 1'b0;  wr_cycle[  963] = 1'b1;  addr_rom[  963]='h00000360;  wr_data_rom[  963]='h000003ea;
    rd_cycle[  964] = 1'b0;  wr_cycle[  964] = 1'b1;  addr_rom[  964]='h0000034c;  wr_data_rom[  964]='h000000c4;
    rd_cycle[  965] = 1'b0;  wr_cycle[  965] = 1'b1;  addr_rom[  965]='h000003b0;  wr_data_rom[  965]='h000001b2;
    rd_cycle[  966] = 1'b0;  wr_cycle[  966] = 1'b1;  addr_rom[  966]='h000003c0;  wr_data_rom[  966]='h00000045;
    rd_cycle[  967] = 1'b0;  wr_cycle[  967] = 1'b1;  addr_rom[  967]='h000001d0;  wr_data_rom[  967]='h00000040;
    rd_cycle[  968] = 1'b0;  wr_cycle[  968] = 1'b1;  addr_rom[  968]='h000002b8;  wr_data_rom[  968]='h000002e0;
    rd_cycle[  969] = 1'b1;  wr_cycle[  969] = 1'b0;  addr_rom[  969]='h000002b8;  wr_data_rom[  969]='h00000000;
    rd_cycle[  970] = 1'b0;  wr_cycle[  970] = 1'b1;  addr_rom[  970]='h00000014;  wr_data_rom[  970]='h0000012f;
    rd_cycle[  971] = 1'b1;  wr_cycle[  971] = 1'b0;  addr_rom[  971]='h00000310;  wr_data_rom[  971]='h00000000;
    rd_cycle[  972] = 1'b0;  wr_cycle[  972] = 1'b1;  addr_rom[  972]='h000002ac;  wr_data_rom[  972]='h000001f1;
    rd_cycle[  973] = 1'b1;  wr_cycle[  973] = 1'b0;  addr_rom[  973]='h000002c4;  wr_data_rom[  973]='h00000000;
    rd_cycle[  974] = 1'b0;  wr_cycle[  974] = 1'b1;  addr_rom[  974]='h000003a4;  wr_data_rom[  974]='h000000fe;
    rd_cycle[  975] = 1'b1;  wr_cycle[  975] = 1'b0;  addr_rom[  975]='h000001e8;  wr_data_rom[  975]='h00000000;
    rd_cycle[  976] = 1'b1;  wr_cycle[  976] = 1'b0;  addr_rom[  976]='h00000084;  wr_data_rom[  976]='h00000000;
    rd_cycle[  977] = 1'b1;  wr_cycle[  977] = 1'b0;  addr_rom[  977]='h000002ac;  wr_data_rom[  977]='h00000000;
    rd_cycle[  978] = 1'b1;  wr_cycle[  978] = 1'b0;  addr_rom[  978]='h00000104;  wr_data_rom[  978]='h00000000;
    rd_cycle[  979] = 1'b1;  wr_cycle[  979] = 1'b0;  addr_rom[  979]='h000001b0;  wr_data_rom[  979]='h00000000;
    rd_cycle[  980] = 1'b1;  wr_cycle[  980] = 1'b0;  addr_rom[  980]='h00000070;  wr_data_rom[  980]='h00000000;
    rd_cycle[  981] = 1'b0;  wr_cycle[  981] = 1'b1;  addr_rom[  981]='h00000008;  wr_data_rom[  981]='h00000237;
    rd_cycle[  982] = 1'b1;  wr_cycle[  982] = 1'b0;  addr_rom[  982]='h000002a8;  wr_data_rom[  982]='h00000000;
    rd_cycle[  983] = 1'b0;  wr_cycle[  983] = 1'b1;  addr_rom[  983]='h00000178;  wr_data_rom[  983]='h0000012f;
    rd_cycle[  984] = 1'b1;  wr_cycle[  984] = 1'b0;  addr_rom[  984]='h000003d8;  wr_data_rom[  984]='h00000000;
    rd_cycle[  985] = 1'b1;  wr_cycle[  985] = 1'b0;  addr_rom[  985]='h00000364;  wr_data_rom[  985]='h00000000;
    rd_cycle[  986] = 1'b0;  wr_cycle[  986] = 1'b1;  addr_rom[  986]='h00000114;  wr_data_rom[  986]='h00000384;
    rd_cycle[  987] = 1'b1;  wr_cycle[  987] = 1'b0;  addr_rom[  987]='h00000340;  wr_data_rom[  987]='h00000000;
    rd_cycle[  988] = 1'b0;  wr_cycle[  988] = 1'b1;  addr_rom[  988]='h000003ac;  wr_data_rom[  988]='h00000088;
    rd_cycle[  989] = 1'b1;  wr_cycle[  989] = 1'b0;  addr_rom[  989]='h00000104;  wr_data_rom[  989]='h00000000;
    rd_cycle[  990] = 1'b1;  wr_cycle[  990] = 1'b0;  addr_rom[  990]='h00000314;  wr_data_rom[  990]='h00000000;
    rd_cycle[  991] = 1'b0;  wr_cycle[  991] = 1'b1;  addr_rom[  991]='h000002a0;  wr_data_rom[  991]='h0000008e;
    rd_cycle[  992] = 1'b0;  wr_cycle[  992] = 1'b1;  addr_rom[  992]='h00000014;  wr_data_rom[  992]='h000001bf;
    rd_cycle[  993] = 1'b1;  wr_cycle[  993] = 1'b0;  addr_rom[  993]='h00000378;  wr_data_rom[  993]='h00000000;
    rd_cycle[  994] = 1'b1;  wr_cycle[  994] = 1'b0;  addr_rom[  994]='h00000178;  wr_data_rom[  994]='h00000000;
    rd_cycle[  995] = 1'b0;  wr_cycle[  995] = 1'b1;  addr_rom[  995]='h00000274;  wr_data_rom[  995]='h000002dc;
    rd_cycle[  996] = 1'b0;  wr_cycle[  996] = 1'b1;  addr_rom[  996]='h00000100;  wr_data_rom[  996]='h00000176;
    rd_cycle[  997] = 1'b0;  wr_cycle[  997] = 1'b1;  addr_rom[  997]='h000003b4;  wr_data_rom[  997]='h00000147;
    rd_cycle[  998] = 1'b0;  wr_cycle[  998] = 1'b1;  addr_rom[  998]='h000000a4;  wr_data_rom[  998]='h00000321;
    rd_cycle[  999] = 1'b1;  wr_cycle[  999] = 1'b0;  addr_rom[  999]='h00000084;  wr_data_rom[  999]='h00000000;
    rd_cycle[ 1000] = 1'b0;  wr_cycle[ 1000] = 1'b1;  addr_rom[ 1000]='h00000260;  wr_data_rom[ 1000]='h000000dd;
    rd_cycle[ 1001] = 1'b1;  wr_cycle[ 1001] = 1'b0;  addr_rom[ 1001]='h000000fc;  wr_data_rom[ 1001]='h00000000;
    rd_cycle[ 1002] = 1'b0;  wr_cycle[ 1002] = 1'b1;  addr_rom[ 1002]='h00000390;  wr_data_rom[ 1002]='h00000050;
    rd_cycle[ 1003] = 1'b0;  wr_cycle[ 1003] = 1'b1;  addr_rom[ 1003]='h000000dc;  wr_data_rom[ 1003]='h000003f1;
    rd_cycle[ 1004] = 1'b1;  wr_cycle[ 1004] = 1'b0;  addr_rom[ 1004]='h00000318;  wr_data_rom[ 1004]='h00000000;
    rd_cycle[ 1005] = 1'b1;  wr_cycle[ 1005] = 1'b0;  addr_rom[ 1005]='h00000224;  wr_data_rom[ 1005]='h00000000;
    rd_cycle[ 1006] = 1'b0;  wr_cycle[ 1006] = 1'b1;  addr_rom[ 1006]='h000001b8;  wr_data_rom[ 1006]='h00000304;
    rd_cycle[ 1007] = 1'b0;  wr_cycle[ 1007] = 1'b1;  addr_rom[ 1007]='h000002d8;  wr_data_rom[ 1007]='h000003ef;
    rd_cycle[ 1008] = 1'b0;  wr_cycle[ 1008] = 1'b1;  addr_rom[ 1008]='h00000394;  wr_data_rom[ 1008]='h000002d6;
    rd_cycle[ 1009] = 1'b0;  wr_cycle[ 1009] = 1'b1;  addr_rom[ 1009]='h0000008c;  wr_data_rom[ 1009]='h00000142;
    rd_cycle[ 1010] = 1'b0;  wr_cycle[ 1010] = 1'b1;  addr_rom[ 1010]='h000000e4;  wr_data_rom[ 1010]='h000003d4;
    rd_cycle[ 1011] = 1'b0;  wr_cycle[ 1011] = 1'b1;  addr_rom[ 1011]='h000001dc;  wr_data_rom[ 1011]='h000002e0;
    rd_cycle[ 1012] = 1'b0;  wr_cycle[ 1012] = 1'b1;  addr_rom[ 1012]='h0000009c;  wr_data_rom[ 1012]='h000002c1;
    rd_cycle[ 1013] = 1'b0;  wr_cycle[ 1013] = 1'b1;  addr_rom[ 1013]='h00000148;  wr_data_rom[ 1013]='h00000367;
    rd_cycle[ 1014] = 1'b0;  wr_cycle[ 1014] = 1'b1;  addr_rom[ 1014]='h0000034c;  wr_data_rom[ 1014]='h00000361;
    rd_cycle[ 1015] = 1'b0;  wr_cycle[ 1015] = 1'b1;  addr_rom[ 1015]='h000002e0;  wr_data_rom[ 1015]='h00000134;
    rd_cycle[ 1016] = 1'b1;  wr_cycle[ 1016] = 1'b0;  addr_rom[ 1016]='h00000168;  wr_data_rom[ 1016]='h00000000;
    rd_cycle[ 1017] = 1'b1;  wr_cycle[ 1017] = 1'b0;  addr_rom[ 1017]='h00000134;  wr_data_rom[ 1017]='h00000000;
    rd_cycle[ 1018] = 1'b1;  wr_cycle[ 1018] = 1'b0;  addr_rom[ 1018]='h00000060;  wr_data_rom[ 1018]='h00000000;
    rd_cycle[ 1019] = 1'b0;  wr_cycle[ 1019] = 1'b1;  addr_rom[ 1019]='h000002d4;  wr_data_rom[ 1019]='h0000005a;
    rd_cycle[ 1020] = 1'b0;  wr_cycle[ 1020] = 1'b1;  addr_rom[ 1020]='h00000388;  wr_data_rom[ 1020]='h00000271;
    rd_cycle[ 1021] = 1'b1;  wr_cycle[ 1021] = 1'b0;  addr_rom[ 1021]='h00000364;  wr_data_rom[ 1021]='h00000000;
    rd_cycle[ 1022] = 1'b1;  wr_cycle[ 1022] = 1'b0;  addr_rom[ 1022]='h00000274;  wr_data_rom[ 1022]='h00000000;
    rd_cycle[ 1023] = 1'b1;  wr_cycle[ 1023] = 1'b0;  addr_rom[ 1023]='h00000064;  wr_data_rom[ 1023]='h00000000;
    // 256 silence cycles
    rd_cycle[ 1024] = 1'b0;  wr_cycle[ 1024] = 1'b0;  addr_rom[ 1024]='h00000000;  wr_data_rom[ 1024]='h00000000;
    rd_cycle[ 1025] = 1'b0;  wr_cycle[ 1025] = 1'b0;  addr_rom[ 1025]='h00000000;  wr_data_rom[ 1025]='h00000000;
    rd_cycle[ 1026] = 1'b0;  wr_cycle[ 1026] = 1'b0;  addr_rom[ 1026]='h00000000;  wr_data_rom[ 1026]='h00000000;
    rd_cycle[ 1027] = 1'b0;  wr_cycle[ 1027] = 1'b0;  addr_rom[ 1027]='h00000000;  wr_data_rom[ 1027]='h00000000;
    rd_cycle[ 1028] = 1'b0;  wr_cycle[ 1028] = 1'b0;  addr_rom[ 1028]='h00000000;  wr_data_rom[ 1028]='h00000000;
    rd_cycle[ 1029] = 1'b0;  wr_cycle[ 1029] = 1'b0;  addr_rom[ 1029]='h00000000;  wr_data_rom[ 1029]='h00000000;
    rd_cycle[ 1030] = 1'b0;  wr_cycle[ 1030] = 1'b0;  addr_rom[ 1030]='h00000000;  wr_data_rom[ 1030]='h00000000;
    rd_cycle[ 1031] = 1'b0;  wr_cycle[ 1031] = 1'b0;  addr_rom[ 1031]='h00000000;  wr_data_rom[ 1031]='h00000000;
    rd_cycle[ 1032] = 1'b0;  wr_cycle[ 1032] = 1'b0;  addr_rom[ 1032]='h00000000;  wr_data_rom[ 1032]='h00000000;
    rd_cycle[ 1033] = 1'b0;  wr_cycle[ 1033] = 1'b0;  addr_rom[ 1033]='h00000000;  wr_data_rom[ 1033]='h00000000;
    rd_cycle[ 1034] = 1'b0;  wr_cycle[ 1034] = 1'b0;  addr_rom[ 1034]='h00000000;  wr_data_rom[ 1034]='h00000000;
    rd_cycle[ 1035] = 1'b0;  wr_cycle[ 1035] = 1'b0;  addr_rom[ 1035]='h00000000;  wr_data_rom[ 1035]='h00000000;
    rd_cycle[ 1036] = 1'b0;  wr_cycle[ 1036] = 1'b0;  addr_rom[ 1036]='h00000000;  wr_data_rom[ 1036]='h00000000;
    rd_cycle[ 1037] = 1'b0;  wr_cycle[ 1037] = 1'b0;  addr_rom[ 1037]='h00000000;  wr_data_rom[ 1037]='h00000000;
    rd_cycle[ 1038] = 1'b0;  wr_cycle[ 1038] = 1'b0;  addr_rom[ 1038]='h00000000;  wr_data_rom[ 1038]='h00000000;
    rd_cycle[ 1039] = 1'b0;  wr_cycle[ 1039] = 1'b0;  addr_rom[ 1039]='h00000000;  wr_data_rom[ 1039]='h00000000;
    rd_cycle[ 1040] = 1'b0;  wr_cycle[ 1040] = 1'b0;  addr_rom[ 1040]='h00000000;  wr_data_rom[ 1040]='h00000000;
    rd_cycle[ 1041] = 1'b0;  wr_cycle[ 1041] = 1'b0;  addr_rom[ 1041]='h00000000;  wr_data_rom[ 1041]='h00000000;
    rd_cycle[ 1042] = 1'b0;  wr_cycle[ 1042] = 1'b0;  addr_rom[ 1042]='h00000000;  wr_data_rom[ 1042]='h00000000;
    rd_cycle[ 1043] = 1'b0;  wr_cycle[ 1043] = 1'b0;  addr_rom[ 1043]='h00000000;  wr_data_rom[ 1043]='h00000000;
    rd_cycle[ 1044] = 1'b0;  wr_cycle[ 1044] = 1'b0;  addr_rom[ 1044]='h00000000;  wr_data_rom[ 1044]='h00000000;
    rd_cycle[ 1045] = 1'b0;  wr_cycle[ 1045] = 1'b0;  addr_rom[ 1045]='h00000000;  wr_data_rom[ 1045]='h00000000;
    rd_cycle[ 1046] = 1'b0;  wr_cycle[ 1046] = 1'b0;  addr_rom[ 1046]='h00000000;  wr_data_rom[ 1046]='h00000000;
    rd_cycle[ 1047] = 1'b0;  wr_cycle[ 1047] = 1'b0;  addr_rom[ 1047]='h00000000;  wr_data_rom[ 1047]='h00000000;
    rd_cycle[ 1048] = 1'b0;  wr_cycle[ 1048] = 1'b0;  addr_rom[ 1048]='h00000000;  wr_data_rom[ 1048]='h00000000;
    rd_cycle[ 1049] = 1'b0;  wr_cycle[ 1049] = 1'b0;  addr_rom[ 1049]='h00000000;  wr_data_rom[ 1049]='h00000000;
    rd_cycle[ 1050] = 1'b0;  wr_cycle[ 1050] = 1'b0;  addr_rom[ 1050]='h00000000;  wr_data_rom[ 1050]='h00000000;
    rd_cycle[ 1051] = 1'b0;  wr_cycle[ 1051] = 1'b0;  addr_rom[ 1051]='h00000000;  wr_data_rom[ 1051]='h00000000;
    rd_cycle[ 1052] = 1'b0;  wr_cycle[ 1052] = 1'b0;  addr_rom[ 1052]='h00000000;  wr_data_rom[ 1052]='h00000000;
    rd_cycle[ 1053] = 1'b0;  wr_cycle[ 1053] = 1'b0;  addr_rom[ 1053]='h00000000;  wr_data_rom[ 1053]='h00000000;
    rd_cycle[ 1054] = 1'b0;  wr_cycle[ 1054] = 1'b0;  addr_rom[ 1054]='h00000000;  wr_data_rom[ 1054]='h00000000;
    rd_cycle[ 1055] = 1'b0;  wr_cycle[ 1055] = 1'b0;  addr_rom[ 1055]='h00000000;  wr_data_rom[ 1055]='h00000000;
    rd_cycle[ 1056] = 1'b0;  wr_cycle[ 1056] = 1'b0;  addr_rom[ 1056]='h00000000;  wr_data_rom[ 1056]='h00000000;
    rd_cycle[ 1057] = 1'b0;  wr_cycle[ 1057] = 1'b0;  addr_rom[ 1057]='h00000000;  wr_data_rom[ 1057]='h00000000;
    rd_cycle[ 1058] = 1'b0;  wr_cycle[ 1058] = 1'b0;  addr_rom[ 1058]='h00000000;  wr_data_rom[ 1058]='h00000000;
    rd_cycle[ 1059] = 1'b0;  wr_cycle[ 1059] = 1'b0;  addr_rom[ 1059]='h00000000;  wr_data_rom[ 1059]='h00000000;
    rd_cycle[ 1060] = 1'b0;  wr_cycle[ 1060] = 1'b0;  addr_rom[ 1060]='h00000000;  wr_data_rom[ 1060]='h00000000;
    rd_cycle[ 1061] = 1'b0;  wr_cycle[ 1061] = 1'b0;  addr_rom[ 1061]='h00000000;  wr_data_rom[ 1061]='h00000000;
    rd_cycle[ 1062] = 1'b0;  wr_cycle[ 1062] = 1'b0;  addr_rom[ 1062]='h00000000;  wr_data_rom[ 1062]='h00000000;
    rd_cycle[ 1063] = 1'b0;  wr_cycle[ 1063] = 1'b0;  addr_rom[ 1063]='h00000000;  wr_data_rom[ 1063]='h00000000;
    rd_cycle[ 1064] = 1'b0;  wr_cycle[ 1064] = 1'b0;  addr_rom[ 1064]='h00000000;  wr_data_rom[ 1064]='h00000000;
    rd_cycle[ 1065] = 1'b0;  wr_cycle[ 1065] = 1'b0;  addr_rom[ 1065]='h00000000;  wr_data_rom[ 1065]='h00000000;
    rd_cycle[ 1066] = 1'b0;  wr_cycle[ 1066] = 1'b0;  addr_rom[ 1066]='h00000000;  wr_data_rom[ 1066]='h00000000;
    rd_cycle[ 1067] = 1'b0;  wr_cycle[ 1067] = 1'b0;  addr_rom[ 1067]='h00000000;  wr_data_rom[ 1067]='h00000000;
    rd_cycle[ 1068] = 1'b0;  wr_cycle[ 1068] = 1'b0;  addr_rom[ 1068]='h00000000;  wr_data_rom[ 1068]='h00000000;
    rd_cycle[ 1069] = 1'b0;  wr_cycle[ 1069] = 1'b0;  addr_rom[ 1069]='h00000000;  wr_data_rom[ 1069]='h00000000;
    rd_cycle[ 1070] = 1'b0;  wr_cycle[ 1070] = 1'b0;  addr_rom[ 1070]='h00000000;  wr_data_rom[ 1070]='h00000000;
    rd_cycle[ 1071] = 1'b0;  wr_cycle[ 1071] = 1'b0;  addr_rom[ 1071]='h00000000;  wr_data_rom[ 1071]='h00000000;
    rd_cycle[ 1072] = 1'b0;  wr_cycle[ 1072] = 1'b0;  addr_rom[ 1072]='h00000000;  wr_data_rom[ 1072]='h00000000;
    rd_cycle[ 1073] = 1'b0;  wr_cycle[ 1073] = 1'b0;  addr_rom[ 1073]='h00000000;  wr_data_rom[ 1073]='h00000000;
    rd_cycle[ 1074] = 1'b0;  wr_cycle[ 1074] = 1'b0;  addr_rom[ 1074]='h00000000;  wr_data_rom[ 1074]='h00000000;
    rd_cycle[ 1075] = 1'b0;  wr_cycle[ 1075] = 1'b0;  addr_rom[ 1075]='h00000000;  wr_data_rom[ 1075]='h00000000;
    rd_cycle[ 1076] = 1'b0;  wr_cycle[ 1076] = 1'b0;  addr_rom[ 1076]='h00000000;  wr_data_rom[ 1076]='h00000000;
    rd_cycle[ 1077] = 1'b0;  wr_cycle[ 1077] = 1'b0;  addr_rom[ 1077]='h00000000;  wr_data_rom[ 1077]='h00000000;
    rd_cycle[ 1078] = 1'b0;  wr_cycle[ 1078] = 1'b0;  addr_rom[ 1078]='h00000000;  wr_data_rom[ 1078]='h00000000;
    rd_cycle[ 1079] = 1'b0;  wr_cycle[ 1079] = 1'b0;  addr_rom[ 1079]='h00000000;  wr_data_rom[ 1079]='h00000000;
    rd_cycle[ 1080] = 1'b0;  wr_cycle[ 1080] = 1'b0;  addr_rom[ 1080]='h00000000;  wr_data_rom[ 1080]='h00000000;
    rd_cycle[ 1081] = 1'b0;  wr_cycle[ 1081] = 1'b0;  addr_rom[ 1081]='h00000000;  wr_data_rom[ 1081]='h00000000;
    rd_cycle[ 1082] = 1'b0;  wr_cycle[ 1082] = 1'b0;  addr_rom[ 1082]='h00000000;  wr_data_rom[ 1082]='h00000000;
    rd_cycle[ 1083] = 1'b0;  wr_cycle[ 1083] = 1'b0;  addr_rom[ 1083]='h00000000;  wr_data_rom[ 1083]='h00000000;
    rd_cycle[ 1084] = 1'b0;  wr_cycle[ 1084] = 1'b0;  addr_rom[ 1084]='h00000000;  wr_data_rom[ 1084]='h00000000;
    rd_cycle[ 1085] = 1'b0;  wr_cycle[ 1085] = 1'b0;  addr_rom[ 1085]='h00000000;  wr_data_rom[ 1085]='h00000000;
    rd_cycle[ 1086] = 1'b0;  wr_cycle[ 1086] = 1'b0;  addr_rom[ 1086]='h00000000;  wr_data_rom[ 1086]='h00000000;
    rd_cycle[ 1087] = 1'b0;  wr_cycle[ 1087] = 1'b0;  addr_rom[ 1087]='h00000000;  wr_data_rom[ 1087]='h00000000;
    rd_cycle[ 1088] = 1'b0;  wr_cycle[ 1088] = 1'b0;  addr_rom[ 1088]='h00000000;  wr_data_rom[ 1088]='h00000000;
    rd_cycle[ 1089] = 1'b0;  wr_cycle[ 1089] = 1'b0;  addr_rom[ 1089]='h00000000;  wr_data_rom[ 1089]='h00000000;
    rd_cycle[ 1090] = 1'b0;  wr_cycle[ 1090] = 1'b0;  addr_rom[ 1090]='h00000000;  wr_data_rom[ 1090]='h00000000;
    rd_cycle[ 1091] = 1'b0;  wr_cycle[ 1091] = 1'b0;  addr_rom[ 1091]='h00000000;  wr_data_rom[ 1091]='h00000000;
    rd_cycle[ 1092] = 1'b0;  wr_cycle[ 1092] = 1'b0;  addr_rom[ 1092]='h00000000;  wr_data_rom[ 1092]='h00000000;
    rd_cycle[ 1093] = 1'b0;  wr_cycle[ 1093] = 1'b0;  addr_rom[ 1093]='h00000000;  wr_data_rom[ 1093]='h00000000;
    rd_cycle[ 1094] = 1'b0;  wr_cycle[ 1094] = 1'b0;  addr_rom[ 1094]='h00000000;  wr_data_rom[ 1094]='h00000000;
    rd_cycle[ 1095] = 1'b0;  wr_cycle[ 1095] = 1'b0;  addr_rom[ 1095]='h00000000;  wr_data_rom[ 1095]='h00000000;
    rd_cycle[ 1096] = 1'b0;  wr_cycle[ 1096] = 1'b0;  addr_rom[ 1096]='h00000000;  wr_data_rom[ 1096]='h00000000;
    rd_cycle[ 1097] = 1'b0;  wr_cycle[ 1097] = 1'b0;  addr_rom[ 1097]='h00000000;  wr_data_rom[ 1097]='h00000000;
    rd_cycle[ 1098] = 1'b0;  wr_cycle[ 1098] = 1'b0;  addr_rom[ 1098]='h00000000;  wr_data_rom[ 1098]='h00000000;
    rd_cycle[ 1099] = 1'b0;  wr_cycle[ 1099] = 1'b0;  addr_rom[ 1099]='h00000000;  wr_data_rom[ 1099]='h00000000;
    rd_cycle[ 1100] = 1'b0;  wr_cycle[ 1100] = 1'b0;  addr_rom[ 1100]='h00000000;  wr_data_rom[ 1100]='h00000000;
    rd_cycle[ 1101] = 1'b0;  wr_cycle[ 1101] = 1'b0;  addr_rom[ 1101]='h00000000;  wr_data_rom[ 1101]='h00000000;
    rd_cycle[ 1102] = 1'b0;  wr_cycle[ 1102] = 1'b0;  addr_rom[ 1102]='h00000000;  wr_data_rom[ 1102]='h00000000;
    rd_cycle[ 1103] = 1'b0;  wr_cycle[ 1103] = 1'b0;  addr_rom[ 1103]='h00000000;  wr_data_rom[ 1103]='h00000000;
    rd_cycle[ 1104] = 1'b0;  wr_cycle[ 1104] = 1'b0;  addr_rom[ 1104]='h00000000;  wr_data_rom[ 1104]='h00000000;
    rd_cycle[ 1105] = 1'b0;  wr_cycle[ 1105] = 1'b0;  addr_rom[ 1105]='h00000000;  wr_data_rom[ 1105]='h00000000;
    rd_cycle[ 1106] = 1'b0;  wr_cycle[ 1106] = 1'b0;  addr_rom[ 1106]='h00000000;  wr_data_rom[ 1106]='h00000000;
    rd_cycle[ 1107] = 1'b0;  wr_cycle[ 1107] = 1'b0;  addr_rom[ 1107]='h00000000;  wr_data_rom[ 1107]='h00000000;
    rd_cycle[ 1108] = 1'b0;  wr_cycle[ 1108] = 1'b0;  addr_rom[ 1108]='h00000000;  wr_data_rom[ 1108]='h00000000;
    rd_cycle[ 1109] = 1'b0;  wr_cycle[ 1109] = 1'b0;  addr_rom[ 1109]='h00000000;  wr_data_rom[ 1109]='h00000000;
    rd_cycle[ 1110] = 1'b0;  wr_cycle[ 1110] = 1'b0;  addr_rom[ 1110]='h00000000;  wr_data_rom[ 1110]='h00000000;
    rd_cycle[ 1111] = 1'b0;  wr_cycle[ 1111] = 1'b0;  addr_rom[ 1111]='h00000000;  wr_data_rom[ 1111]='h00000000;
    rd_cycle[ 1112] = 1'b0;  wr_cycle[ 1112] = 1'b0;  addr_rom[ 1112]='h00000000;  wr_data_rom[ 1112]='h00000000;
    rd_cycle[ 1113] = 1'b0;  wr_cycle[ 1113] = 1'b0;  addr_rom[ 1113]='h00000000;  wr_data_rom[ 1113]='h00000000;
    rd_cycle[ 1114] = 1'b0;  wr_cycle[ 1114] = 1'b0;  addr_rom[ 1114]='h00000000;  wr_data_rom[ 1114]='h00000000;
    rd_cycle[ 1115] = 1'b0;  wr_cycle[ 1115] = 1'b0;  addr_rom[ 1115]='h00000000;  wr_data_rom[ 1115]='h00000000;
    rd_cycle[ 1116] = 1'b0;  wr_cycle[ 1116] = 1'b0;  addr_rom[ 1116]='h00000000;  wr_data_rom[ 1116]='h00000000;
    rd_cycle[ 1117] = 1'b0;  wr_cycle[ 1117] = 1'b0;  addr_rom[ 1117]='h00000000;  wr_data_rom[ 1117]='h00000000;
    rd_cycle[ 1118] = 1'b0;  wr_cycle[ 1118] = 1'b0;  addr_rom[ 1118]='h00000000;  wr_data_rom[ 1118]='h00000000;
    rd_cycle[ 1119] = 1'b0;  wr_cycle[ 1119] = 1'b0;  addr_rom[ 1119]='h00000000;  wr_data_rom[ 1119]='h00000000;
    rd_cycle[ 1120] = 1'b0;  wr_cycle[ 1120] = 1'b0;  addr_rom[ 1120]='h00000000;  wr_data_rom[ 1120]='h00000000;
    rd_cycle[ 1121] = 1'b0;  wr_cycle[ 1121] = 1'b0;  addr_rom[ 1121]='h00000000;  wr_data_rom[ 1121]='h00000000;
    rd_cycle[ 1122] = 1'b0;  wr_cycle[ 1122] = 1'b0;  addr_rom[ 1122]='h00000000;  wr_data_rom[ 1122]='h00000000;
    rd_cycle[ 1123] = 1'b0;  wr_cycle[ 1123] = 1'b0;  addr_rom[ 1123]='h00000000;  wr_data_rom[ 1123]='h00000000;
    rd_cycle[ 1124] = 1'b0;  wr_cycle[ 1124] = 1'b0;  addr_rom[ 1124]='h00000000;  wr_data_rom[ 1124]='h00000000;
    rd_cycle[ 1125] = 1'b0;  wr_cycle[ 1125] = 1'b0;  addr_rom[ 1125]='h00000000;  wr_data_rom[ 1125]='h00000000;
    rd_cycle[ 1126] = 1'b0;  wr_cycle[ 1126] = 1'b0;  addr_rom[ 1126]='h00000000;  wr_data_rom[ 1126]='h00000000;
    rd_cycle[ 1127] = 1'b0;  wr_cycle[ 1127] = 1'b0;  addr_rom[ 1127]='h00000000;  wr_data_rom[ 1127]='h00000000;
    rd_cycle[ 1128] = 1'b0;  wr_cycle[ 1128] = 1'b0;  addr_rom[ 1128]='h00000000;  wr_data_rom[ 1128]='h00000000;
    rd_cycle[ 1129] = 1'b0;  wr_cycle[ 1129] = 1'b0;  addr_rom[ 1129]='h00000000;  wr_data_rom[ 1129]='h00000000;
    rd_cycle[ 1130] = 1'b0;  wr_cycle[ 1130] = 1'b0;  addr_rom[ 1130]='h00000000;  wr_data_rom[ 1130]='h00000000;
    rd_cycle[ 1131] = 1'b0;  wr_cycle[ 1131] = 1'b0;  addr_rom[ 1131]='h00000000;  wr_data_rom[ 1131]='h00000000;
    rd_cycle[ 1132] = 1'b0;  wr_cycle[ 1132] = 1'b0;  addr_rom[ 1132]='h00000000;  wr_data_rom[ 1132]='h00000000;
    rd_cycle[ 1133] = 1'b0;  wr_cycle[ 1133] = 1'b0;  addr_rom[ 1133]='h00000000;  wr_data_rom[ 1133]='h00000000;
    rd_cycle[ 1134] = 1'b0;  wr_cycle[ 1134] = 1'b0;  addr_rom[ 1134]='h00000000;  wr_data_rom[ 1134]='h00000000;
    rd_cycle[ 1135] = 1'b0;  wr_cycle[ 1135] = 1'b0;  addr_rom[ 1135]='h00000000;  wr_data_rom[ 1135]='h00000000;
    rd_cycle[ 1136] = 1'b0;  wr_cycle[ 1136] = 1'b0;  addr_rom[ 1136]='h00000000;  wr_data_rom[ 1136]='h00000000;
    rd_cycle[ 1137] = 1'b0;  wr_cycle[ 1137] = 1'b0;  addr_rom[ 1137]='h00000000;  wr_data_rom[ 1137]='h00000000;
    rd_cycle[ 1138] = 1'b0;  wr_cycle[ 1138] = 1'b0;  addr_rom[ 1138]='h00000000;  wr_data_rom[ 1138]='h00000000;
    rd_cycle[ 1139] = 1'b0;  wr_cycle[ 1139] = 1'b0;  addr_rom[ 1139]='h00000000;  wr_data_rom[ 1139]='h00000000;
    rd_cycle[ 1140] = 1'b0;  wr_cycle[ 1140] = 1'b0;  addr_rom[ 1140]='h00000000;  wr_data_rom[ 1140]='h00000000;
    rd_cycle[ 1141] = 1'b0;  wr_cycle[ 1141] = 1'b0;  addr_rom[ 1141]='h00000000;  wr_data_rom[ 1141]='h00000000;
    rd_cycle[ 1142] = 1'b0;  wr_cycle[ 1142] = 1'b0;  addr_rom[ 1142]='h00000000;  wr_data_rom[ 1142]='h00000000;
    rd_cycle[ 1143] = 1'b0;  wr_cycle[ 1143] = 1'b0;  addr_rom[ 1143]='h00000000;  wr_data_rom[ 1143]='h00000000;
    rd_cycle[ 1144] = 1'b0;  wr_cycle[ 1144] = 1'b0;  addr_rom[ 1144]='h00000000;  wr_data_rom[ 1144]='h00000000;
    rd_cycle[ 1145] = 1'b0;  wr_cycle[ 1145] = 1'b0;  addr_rom[ 1145]='h00000000;  wr_data_rom[ 1145]='h00000000;
    rd_cycle[ 1146] = 1'b0;  wr_cycle[ 1146] = 1'b0;  addr_rom[ 1146]='h00000000;  wr_data_rom[ 1146]='h00000000;
    rd_cycle[ 1147] = 1'b0;  wr_cycle[ 1147] = 1'b0;  addr_rom[ 1147]='h00000000;  wr_data_rom[ 1147]='h00000000;
    rd_cycle[ 1148] = 1'b0;  wr_cycle[ 1148] = 1'b0;  addr_rom[ 1148]='h00000000;  wr_data_rom[ 1148]='h00000000;
    rd_cycle[ 1149] = 1'b0;  wr_cycle[ 1149] = 1'b0;  addr_rom[ 1149]='h00000000;  wr_data_rom[ 1149]='h00000000;
    rd_cycle[ 1150] = 1'b0;  wr_cycle[ 1150] = 1'b0;  addr_rom[ 1150]='h00000000;  wr_data_rom[ 1150]='h00000000;
    rd_cycle[ 1151] = 1'b0;  wr_cycle[ 1151] = 1'b0;  addr_rom[ 1151]='h00000000;  wr_data_rom[ 1151]='h00000000;
    rd_cycle[ 1152] = 1'b0;  wr_cycle[ 1152] = 1'b0;  addr_rom[ 1152]='h00000000;  wr_data_rom[ 1152]='h00000000;
    rd_cycle[ 1153] = 1'b0;  wr_cycle[ 1153] = 1'b0;  addr_rom[ 1153]='h00000000;  wr_data_rom[ 1153]='h00000000;
    rd_cycle[ 1154] = 1'b0;  wr_cycle[ 1154] = 1'b0;  addr_rom[ 1154]='h00000000;  wr_data_rom[ 1154]='h00000000;
    rd_cycle[ 1155] = 1'b0;  wr_cycle[ 1155] = 1'b0;  addr_rom[ 1155]='h00000000;  wr_data_rom[ 1155]='h00000000;
    rd_cycle[ 1156] = 1'b0;  wr_cycle[ 1156] = 1'b0;  addr_rom[ 1156]='h00000000;  wr_data_rom[ 1156]='h00000000;
    rd_cycle[ 1157] = 1'b0;  wr_cycle[ 1157] = 1'b0;  addr_rom[ 1157]='h00000000;  wr_data_rom[ 1157]='h00000000;
    rd_cycle[ 1158] = 1'b0;  wr_cycle[ 1158] = 1'b0;  addr_rom[ 1158]='h00000000;  wr_data_rom[ 1158]='h00000000;
    rd_cycle[ 1159] = 1'b0;  wr_cycle[ 1159] = 1'b0;  addr_rom[ 1159]='h00000000;  wr_data_rom[ 1159]='h00000000;
    rd_cycle[ 1160] = 1'b0;  wr_cycle[ 1160] = 1'b0;  addr_rom[ 1160]='h00000000;  wr_data_rom[ 1160]='h00000000;
    rd_cycle[ 1161] = 1'b0;  wr_cycle[ 1161] = 1'b0;  addr_rom[ 1161]='h00000000;  wr_data_rom[ 1161]='h00000000;
    rd_cycle[ 1162] = 1'b0;  wr_cycle[ 1162] = 1'b0;  addr_rom[ 1162]='h00000000;  wr_data_rom[ 1162]='h00000000;
    rd_cycle[ 1163] = 1'b0;  wr_cycle[ 1163] = 1'b0;  addr_rom[ 1163]='h00000000;  wr_data_rom[ 1163]='h00000000;
    rd_cycle[ 1164] = 1'b0;  wr_cycle[ 1164] = 1'b0;  addr_rom[ 1164]='h00000000;  wr_data_rom[ 1164]='h00000000;
    rd_cycle[ 1165] = 1'b0;  wr_cycle[ 1165] = 1'b0;  addr_rom[ 1165]='h00000000;  wr_data_rom[ 1165]='h00000000;
    rd_cycle[ 1166] = 1'b0;  wr_cycle[ 1166] = 1'b0;  addr_rom[ 1166]='h00000000;  wr_data_rom[ 1166]='h00000000;
    rd_cycle[ 1167] = 1'b0;  wr_cycle[ 1167] = 1'b0;  addr_rom[ 1167]='h00000000;  wr_data_rom[ 1167]='h00000000;
    rd_cycle[ 1168] = 1'b0;  wr_cycle[ 1168] = 1'b0;  addr_rom[ 1168]='h00000000;  wr_data_rom[ 1168]='h00000000;
    rd_cycle[ 1169] = 1'b0;  wr_cycle[ 1169] = 1'b0;  addr_rom[ 1169]='h00000000;  wr_data_rom[ 1169]='h00000000;
    rd_cycle[ 1170] = 1'b0;  wr_cycle[ 1170] = 1'b0;  addr_rom[ 1170]='h00000000;  wr_data_rom[ 1170]='h00000000;
    rd_cycle[ 1171] = 1'b0;  wr_cycle[ 1171] = 1'b0;  addr_rom[ 1171]='h00000000;  wr_data_rom[ 1171]='h00000000;
    rd_cycle[ 1172] = 1'b0;  wr_cycle[ 1172] = 1'b0;  addr_rom[ 1172]='h00000000;  wr_data_rom[ 1172]='h00000000;
    rd_cycle[ 1173] = 1'b0;  wr_cycle[ 1173] = 1'b0;  addr_rom[ 1173]='h00000000;  wr_data_rom[ 1173]='h00000000;
    rd_cycle[ 1174] = 1'b0;  wr_cycle[ 1174] = 1'b0;  addr_rom[ 1174]='h00000000;  wr_data_rom[ 1174]='h00000000;
    rd_cycle[ 1175] = 1'b0;  wr_cycle[ 1175] = 1'b0;  addr_rom[ 1175]='h00000000;  wr_data_rom[ 1175]='h00000000;
    rd_cycle[ 1176] = 1'b0;  wr_cycle[ 1176] = 1'b0;  addr_rom[ 1176]='h00000000;  wr_data_rom[ 1176]='h00000000;
    rd_cycle[ 1177] = 1'b0;  wr_cycle[ 1177] = 1'b0;  addr_rom[ 1177]='h00000000;  wr_data_rom[ 1177]='h00000000;
    rd_cycle[ 1178] = 1'b0;  wr_cycle[ 1178] = 1'b0;  addr_rom[ 1178]='h00000000;  wr_data_rom[ 1178]='h00000000;
    rd_cycle[ 1179] = 1'b0;  wr_cycle[ 1179] = 1'b0;  addr_rom[ 1179]='h00000000;  wr_data_rom[ 1179]='h00000000;
    rd_cycle[ 1180] = 1'b0;  wr_cycle[ 1180] = 1'b0;  addr_rom[ 1180]='h00000000;  wr_data_rom[ 1180]='h00000000;
    rd_cycle[ 1181] = 1'b0;  wr_cycle[ 1181] = 1'b0;  addr_rom[ 1181]='h00000000;  wr_data_rom[ 1181]='h00000000;
    rd_cycle[ 1182] = 1'b0;  wr_cycle[ 1182] = 1'b0;  addr_rom[ 1182]='h00000000;  wr_data_rom[ 1182]='h00000000;
    rd_cycle[ 1183] = 1'b0;  wr_cycle[ 1183] = 1'b0;  addr_rom[ 1183]='h00000000;  wr_data_rom[ 1183]='h00000000;
    rd_cycle[ 1184] = 1'b0;  wr_cycle[ 1184] = 1'b0;  addr_rom[ 1184]='h00000000;  wr_data_rom[ 1184]='h00000000;
    rd_cycle[ 1185] = 1'b0;  wr_cycle[ 1185] = 1'b0;  addr_rom[ 1185]='h00000000;  wr_data_rom[ 1185]='h00000000;
    rd_cycle[ 1186] = 1'b0;  wr_cycle[ 1186] = 1'b0;  addr_rom[ 1186]='h00000000;  wr_data_rom[ 1186]='h00000000;
    rd_cycle[ 1187] = 1'b0;  wr_cycle[ 1187] = 1'b0;  addr_rom[ 1187]='h00000000;  wr_data_rom[ 1187]='h00000000;
    rd_cycle[ 1188] = 1'b0;  wr_cycle[ 1188] = 1'b0;  addr_rom[ 1188]='h00000000;  wr_data_rom[ 1188]='h00000000;
    rd_cycle[ 1189] = 1'b0;  wr_cycle[ 1189] = 1'b0;  addr_rom[ 1189]='h00000000;  wr_data_rom[ 1189]='h00000000;
    rd_cycle[ 1190] = 1'b0;  wr_cycle[ 1190] = 1'b0;  addr_rom[ 1190]='h00000000;  wr_data_rom[ 1190]='h00000000;
    rd_cycle[ 1191] = 1'b0;  wr_cycle[ 1191] = 1'b0;  addr_rom[ 1191]='h00000000;  wr_data_rom[ 1191]='h00000000;
    rd_cycle[ 1192] = 1'b0;  wr_cycle[ 1192] = 1'b0;  addr_rom[ 1192]='h00000000;  wr_data_rom[ 1192]='h00000000;
    rd_cycle[ 1193] = 1'b0;  wr_cycle[ 1193] = 1'b0;  addr_rom[ 1193]='h00000000;  wr_data_rom[ 1193]='h00000000;
    rd_cycle[ 1194] = 1'b0;  wr_cycle[ 1194] = 1'b0;  addr_rom[ 1194]='h00000000;  wr_data_rom[ 1194]='h00000000;
    rd_cycle[ 1195] = 1'b0;  wr_cycle[ 1195] = 1'b0;  addr_rom[ 1195]='h00000000;  wr_data_rom[ 1195]='h00000000;
    rd_cycle[ 1196] = 1'b0;  wr_cycle[ 1196] = 1'b0;  addr_rom[ 1196]='h00000000;  wr_data_rom[ 1196]='h00000000;
    rd_cycle[ 1197] = 1'b0;  wr_cycle[ 1197] = 1'b0;  addr_rom[ 1197]='h00000000;  wr_data_rom[ 1197]='h00000000;
    rd_cycle[ 1198] = 1'b0;  wr_cycle[ 1198] = 1'b0;  addr_rom[ 1198]='h00000000;  wr_data_rom[ 1198]='h00000000;
    rd_cycle[ 1199] = 1'b0;  wr_cycle[ 1199] = 1'b0;  addr_rom[ 1199]='h00000000;  wr_data_rom[ 1199]='h00000000;
    rd_cycle[ 1200] = 1'b0;  wr_cycle[ 1200] = 1'b0;  addr_rom[ 1200]='h00000000;  wr_data_rom[ 1200]='h00000000;
    rd_cycle[ 1201] = 1'b0;  wr_cycle[ 1201] = 1'b0;  addr_rom[ 1201]='h00000000;  wr_data_rom[ 1201]='h00000000;
    rd_cycle[ 1202] = 1'b0;  wr_cycle[ 1202] = 1'b0;  addr_rom[ 1202]='h00000000;  wr_data_rom[ 1202]='h00000000;
    rd_cycle[ 1203] = 1'b0;  wr_cycle[ 1203] = 1'b0;  addr_rom[ 1203]='h00000000;  wr_data_rom[ 1203]='h00000000;
    rd_cycle[ 1204] = 1'b0;  wr_cycle[ 1204] = 1'b0;  addr_rom[ 1204]='h00000000;  wr_data_rom[ 1204]='h00000000;
    rd_cycle[ 1205] = 1'b0;  wr_cycle[ 1205] = 1'b0;  addr_rom[ 1205]='h00000000;  wr_data_rom[ 1205]='h00000000;
    rd_cycle[ 1206] = 1'b0;  wr_cycle[ 1206] = 1'b0;  addr_rom[ 1206]='h00000000;  wr_data_rom[ 1206]='h00000000;
    rd_cycle[ 1207] = 1'b0;  wr_cycle[ 1207] = 1'b0;  addr_rom[ 1207]='h00000000;  wr_data_rom[ 1207]='h00000000;
    rd_cycle[ 1208] = 1'b0;  wr_cycle[ 1208] = 1'b0;  addr_rom[ 1208]='h00000000;  wr_data_rom[ 1208]='h00000000;
    rd_cycle[ 1209] = 1'b0;  wr_cycle[ 1209] = 1'b0;  addr_rom[ 1209]='h00000000;  wr_data_rom[ 1209]='h00000000;
    rd_cycle[ 1210] = 1'b0;  wr_cycle[ 1210] = 1'b0;  addr_rom[ 1210]='h00000000;  wr_data_rom[ 1210]='h00000000;
    rd_cycle[ 1211] = 1'b0;  wr_cycle[ 1211] = 1'b0;  addr_rom[ 1211]='h00000000;  wr_data_rom[ 1211]='h00000000;
    rd_cycle[ 1212] = 1'b0;  wr_cycle[ 1212] = 1'b0;  addr_rom[ 1212]='h00000000;  wr_data_rom[ 1212]='h00000000;
    rd_cycle[ 1213] = 1'b0;  wr_cycle[ 1213] = 1'b0;  addr_rom[ 1213]='h00000000;  wr_data_rom[ 1213]='h00000000;
    rd_cycle[ 1214] = 1'b0;  wr_cycle[ 1214] = 1'b0;  addr_rom[ 1214]='h00000000;  wr_data_rom[ 1214]='h00000000;
    rd_cycle[ 1215] = 1'b0;  wr_cycle[ 1215] = 1'b0;  addr_rom[ 1215]='h00000000;  wr_data_rom[ 1215]='h00000000;
    rd_cycle[ 1216] = 1'b0;  wr_cycle[ 1216] = 1'b0;  addr_rom[ 1216]='h00000000;  wr_data_rom[ 1216]='h00000000;
    rd_cycle[ 1217] = 1'b0;  wr_cycle[ 1217] = 1'b0;  addr_rom[ 1217]='h00000000;  wr_data_rom[ 1217]='h00000000;
    rd_cycle[ 1218] = 1'b0;  wr_cycle[ 1218] = 1'b0;  addr_rom[ 1218]='h00000000;  wr_data_rom[ 1218]='h00000000;
    rd_cycle[ 1219] = 1'b0;  wr_cycle[ 1219] = 1'b0;  addr_rom[ 1219]='h00000000;  wr_data_rom[ 1219]='h00000000;
    rd_cycle[ 1220] = 1'b0;  wr_cycle[ 1220] = 1'b0;  addr_rom[ 1220]='h00000000;  wr_data_rom[ 1220]='h00000000;
    rd_cycle[ 1221] = 1'b0;  wr_cycle[ 1221] = 1'b0;  addr_rom[ 1221]='h00000000;  wr_data_rom[ 1221]='h00000000;
    rd_cycle[ 1222] = 1'b0;  wr_cycle[ 1222] = 1'b0;  addr_rom[ 1222]='h00000000;  wr_data_rom[ 1222]='h00000000;
    rd_cycle[ 1223] = 1'b0;  wr_cycle[ 1223] = 1'b0;  addr_rom[ 1223]='h00000000;  wr_data_rom[ 1223]='h00000000;
    rd_cycle[ 1224] = 1'b0;  wr_cycle[ 1224] = 1'b0;  addr_rom[ 1224]='h00000000;  wr_data_rom[ 1224]='h00000000;
    rd_cycle[ 1225] = 1'b0;  wr_cycle[ 1225] = 1'b0;  addr_rom[ 1225]='h00000000;  wr_data_rom[ 1225]='h00000000;
    rd_cycle[ 1226] = 1'b0;  wr_cycle[ 1226] = 1'b0;  addr_rom[ 1226]='h00000000;  wr_data_rom[ 1226]='h00000000;
    rd_cycle[ 1227] = 1'b0;  wr_cycle[ 1227] = 1'b0;  addr_rom[ 1227]='h00000000;  wr_data_rom[ 1227]='h00000000;
    rd_cycle[ 1228] = 1'b0;  wr_cycle[ 1228] = 1'b0;  addr_rom[ 1228]='h00000000;  wr_data_rom[ 1228]='h00000000;
    rd_cycle[ 1229] = 1'b0;  wr_cycle[ 1229] = 1'b0;  addr_rom[ 1229]='h00000000;  wr_data_rom[ 1229]='h00000000;
    rd_cycle[ 1230] = 1'b0;  wr_cycle[ 1230] = 1'b0;  addr_rom[ 1230]='h00000000;  wr_data_rom[ 1230]='h00000000;
    rd_cycle[ 1231] = 1'b0;  wr_cycle[ 1231] = 1'b0;  addr_rom[ 1231]='h00000000;  wr_data_rom[ 1231]='h00000000;
    rd_cycle[ 1232] = 1'b0;  wr_cycle[ 1232] = 1'b0;  addr_rom[ 1232]='h00000000;  wr_data_rom[ 1232]='h00000000;
    rd_cycle[ 1233] = 1'b0;  wr_cycle[ 1233] = 1'b0;  addr_rom[ 1233]='h00000000;  wr_data_rom[ 1233]='h00000000;
    rd_cycle[ 1234] = 1'b0;  wr_cycle[ 1234] = 1'b0;  addr_rom[ 1234]='h00000000;  wr_data_rom[ 1234]='h00000000;
    rd_cycle[ 1235] = 1'b0;  wr_cycle[ 1235] = 1'b0;  addr_rom[ 1235]='h00000000;  wr_data_rom[ 1235]='h00000000;
    rd_cycle[ 1236] = 1'b0;  wr_cycle[ 1236] = 1'b0;  addr_rom[ 1236]='h00000000;  wr_data_rom[ 1236]='h00000000;
    rd_cycle[ 1237] = 1'b0;  wr_cycle[ 1237] = 1'b0;  addr_rom[ 1237]='h00000000;  wr_data_rom[ 1237]='h00000000;
    rd_cycle[ 1238] = 1'b0;  wr_cycle[ 1238] = 1'b0;  addr_rom[ 1238]='h00000000;  wr_data_rom[ 1238]='h00000000;
    rd_cycle[ 1239] = 1'b0;  wr_cycle[ 1239] = 1'b0;  addr_rom[ 1239]='h00000000;  wr_data_rom[ 1239]='h00000000;
    rd_cycle[ 1240] = 1'b0;  wr_cycle[ 1240] = 1'b0;  addr_rom[ 1240]='h00000000;  wr_data_rom[ 1240]='h00000000;
    rd_cycle[ 1241] = 1'b0;  wr_cycle[ 1241] = 1'b0;  addr_rom[ 1241]='h00000000;  wr_data_rom[ 1241]='h00000000;
    rd_cycle[ 1242] = 1'b0;  wr_cycle[ 1242] = 1'b0;  addr_rom[ 1242]='h00000000;  wr_data_rom[ 1242]='h00000000;
    rd_cycle[ 1243] = 1'b0;  wr_cycle[ 1243] = 1'b0;  addr_rom[ 1243]='h00000000;  wr_data_rom[ 1243]='h00000000;
    rd_cycle[ 1244] = 1'b0;  wr_cycle[ 1244] = 1'b0;  addr_rom[ 1244]='h00000000;  wr_data_rom[ 1244]='h00000000;
    rd_cycle[ 1245] = 1'b0;  wr_cycle[ 1245] = 1'b0;  addr_rom[ 1245]='h00000000;  wr_data_rom[ 1245]='h00000000;
    rd_cycle[ 1246] = 1'b0;  wr_cycle[ 1246] = 1'b0;  addr_rom[ 1246]='h00000000;  wr_data_rom[ 1246]='h00000000;
    rd_cycle[ 1247] = 1'b0;  wr_cycle[ 1247] = 1'b0;  addr_rom[ 1247]='h00000000;  wr_data_rom[ 1247]='h00000000;
    rd_cycle[ 1248] = 1'b0;  wr_cycle[ 1248] = 1'b0;  addr_rom[ 1248]='h00000000;  wr_data_rom[ 1248]='h00000000;
    rd_cycle[ 1249] = 1'b0;  wr_cycle[ 1249] = 1'b0;  addr_rom[ 1249]='h00000000;  wr_data_rom[ 1249]='h00000000;
    rd_cycle[ 1250] = 1'b0;  wr_cycle[ 1250] = 1'b0;  addr_rom[ 1250]='h00000000;  wr_data_rom[ 1250]='h00000000;
    rd_cycle[ 1251] = 1'b0;  wr_cycle[ 1251] = 1'b0;  addr_rom[ 1251]='h00000000;  wr_data_rom[ 1251]='h00000000;
    rd_cycle[ 1252] = 1'b0;  wr_cycle[ 1252] = 1'b0;  addr_rom[ 1252]='h00000000;  wr_data_rom[ 1252]='h00000000;
    rd_cycle[ 1253] = 1'b0;  wr_cycle[ 1253] = 1'b0;  addr_rom[ 1253]='h00000000;  wr_data_rom[ 1253]='h00000000;
    rd_cycle[ 1254] = 1'b0;  wr_cycle[ 1254] = 1'b0;  addr_rom[ 1254]='h00000000;  wr_data_rom[ 1254]='h00000000;
    rd_cycle[ 1255] = 1'b0;  wr_cycle[ 1255] = 1'b0;  addr_rom[ 1255]='h00000000;  wr_data_rom[ 1255]='h00000000;
    rd_cycle[ 1256] = 1'b0;  wr_cycle[ 1256] = 1'b0;  addr_rom[ 1256]='h00000000;  wr_data_rom[ 1256]='h00000000;
    rd_cycle[ 1257] = 1'b0;  wr_cycle[ 1257] = 1'b0;  addr_rom[ 1257]='h00000000;  wr_data_rom[ 1257]='h00000000;
    rd_cycle[ 1258] = 1'b0;  wr_cycle[ 1258] = 1'b0;  addr_rom[ 1258]='h00000000;  wr_data_rom[ 1258]='h00000000;
    rd_cycle[ 1259] = 1'b0;  wr_cycle[ 1259] = 1'b0;  addr_rom[ 1259]='h00000000;  wr_data_rom[ 1259]='h00000000;
    rd_cycle[ 1260] = 1'b0;  wr_cycle[ 1260] = 1'b0;  addr_rom[ 1260]='h00000000;  wr_data_rom[ 1260]='h00000000;
    rd_cycle[ 1261] = 1'b0;  wr_cycle[ 1261] = 1'b0;  addr_rom[ 1261]='h00000000;  wr_data_rom[ 1261]='h00000000;
    rd_cycle[ 1262] = 1'b0;  wr_cycle[ 1262] = 1'b0;  addr_rom[ 1262]='h00000000;  wr_data_rom[ 1262]='h00000000;
    rd_cycle[ 1263] = 1'b0;  wr_cycle[ 1263] = 1'b0;  addr_rom[ 1263]='h00000000;  wr_data_rom[ 1263]='h00000000;
    rd_cycle[ 1264] = 1'b0;  wr_cycle[ 1264] = 1'b0;  addr_rom[ 1264]='h00000000;  wr_data_rom[ 1264]='h00000000;
    rd_cycle[ 1265] = 1'b0;  wr_cycle[ 1265] = 1'b0;  addr_rom[ 1265]='h00000000;  wr_data_rom[ 1265]='h00000000;
    rd_cycle[ 1266] = 1'b0;  wr_cycle[ 1266] = 1'b0;  addr_rom[ 1266]='h00000000;  wr_data_rom[ 1266]='h00000000;
    rd_cycle[ 1267] = 1'b0;  wr_cycle[ 1267] = 1'b0;  addr_rom[ 1267]='h00000000;  wr_data_rom[ 1267]='h00000000;
    rd_cycle[ 1268] = 1'b0;  wr_cycle[ 1268] = 1'b0;  addr_rom[ 1268]='h00000000;  wr_data_rom[ 1268]='h00000000;
    rd_cycle[ 1269] = 1'b0;  wr_cycle[ 1269] = 1'b0;  addr_rom[ 1269]='h00000000;  wr_data_rom[ 1269]='h00000000;
    rd_cycle[ 1270] = 1'b0;  wr_cycle[ 1270] = 1'b0;  addr_rom[ 1270]='h00000000;  wr_data_rom[ 1270]='h00000000;
    rd_cycle[ 1271] = 1'b0;  wr_cycle[ 1271] = 1'b0;  addr_rom[ 1271]='h00000000;  wr_data_rom[ 1271]='h00000000;
    rd_cycle[ 1272] = 1'b0;  wr_cycle[ 1272] = 1'b0;  addr_rom[ 1272]='h00000000;  wr_data_rom[ 1272]='h00000000;
    rd_cycle[ 1273] = 1'b0;  wr_cycle[ 1273] = 1'b0;  addr_rom[ 1273]='h00000000;  wr_data_rom[ 1273]='h00000000;
    rd_cycle[ 1274] = 1'b0;  wr_cycle[ 1274] = 1'b0;  addr_rom[ 1274]='h00000000;  wr_data_rom[ 1274]='h00000000;
    rd_cycle[ 1275] = 1'b0;  wr_cycle[ 1275] = 1'b0;  addr_rom[ 1275]='h00000000;  wr_data_rom[ 1275]='h00000000;
    rd_cycle[ 1276] = 1'b0;  wr_cycle[ 1276] = 1'b0;  addr_rom[ 1276]='h00000000;  wr_data_rom[ 1276]='h00000000;
    rd_cycle[ 1277] = 1'b0;  wr_cycle[ 1277] = 1'b0;  addr_rom[ 1277]='h00000000;  wr_data_rom[ 1277]='h00000000;
    rd_cycle[ 1278] = 1'b0;  wr_cycle[ 1278] = 1'b0;  addr_rom[ 1278]='h00000000;  wr_data_rom[ 1278]='h00000000;
    rd_cycle[ 1279] = 1'b0;  wr_cycle[ 1279] = 1'b0;  addr_rom[ 1279]='h00000000;  wr_data_rom[ 1279]='h00000000;
    // 256 sequence read cycles
    rd_cycle[ 1280] = 1'b1;  wr_cycle[ 1280] = 1'b0;  addr_rom[ 1280]='h00000000;  wr_data_rom[ 1280]='h00000000;
    rd_cycle[ 1281] = 1'b1;  wr_cycle[ 1281] = 1'b0;  addr_rom[ 1281]='h00000004;  wr_data_rom[ 1281]='h00000000;
    rd_cycle[ 1282] = 1'b1;  wr_cycle[ 1282] = 1'b0;  addr_rom[ 1282]='h00000008;  wr_data_rom[ 1282]='h00000000;
    rd_cycle[ 1283] = 1'b1;  wr_cycle[ 1283] = 1'b0;  addr_rom[ 1283]='h0000000c;  wr_data_rom[ 1283]='h00000000;
    rd_cycle[ 1284] = 1'b1;  wr_cycle[ 1284] = 1'b0;  addr_rom[ 1284]='h00000010;  wr_data_rom[ 1284]='h00000000;
    rd_cycle[ 1285] = 1'b1;  wr_cycle[ 1285] = 1'b0;  addr_rom[ 1285]='h00000014;  wr_data_rom[ 1285]='h00000000;
    rd_cycle[ 1286] = 1'b1;  wr_cycle[ 1286] = 1'b0;  addr_rom[ 1286]='h00000018;  wr_data_rom[ 1286]='h00000000;
    rd_cycle[ 1287] = 1'b1;  wr_cycle[ 1287] = 1'b0;  addr_rom[ 1287]='h0000001c;  wr_data_rom[ 1287]='h00000000;
    rd_cycle[ 1288] = 1'b1;  wr_cycle[ 1288] = 1'b0;  addr_rom[ 1288]='h00000020;  wr_data_rom[ 1288]='h00000000;
    rd_cycle[ 1289] = 1'b1;  wr_cycle[ 1289] = 1'b0;  addr_rom[ 1289]='h00000024;  wr_data_rom[ 1289]='h00000000;
    rd_cycle[ 1290] = 1'b1;  wr_cycle[ 1290] = 1'b0;  addr_rom[ 1290]='h00000028;  wr_data_rom[ 1290]='h00000000;
    rd_cycle[ 1291] = 1'b1;  wr_cycle[ 1291] = 1'b0;  addr_rom[ 1291]='h0000002c;  wr_data_rom[ 1291]='h00000000;
    rd_cycle[ 1292] = 1'b1;  wr_cycle[ 1292] = 1'b0;  addr_rom[ 1292]='h00000030;  wr_data_rom[ 1292]='h00000000;
    rd_cycle[ 1293] = 1'b1;  wr_cycle[ 1293] = 1'b0;  addr_rom[ 1293]='h00000034;  wr_data_rom[ 1293]='h00000000;
    rd_cycle[ 1294] = 1'b1;  wr_cycle[ 1294] = 1'b0;  addr_rom[ 1294]='h00000038;  wr_data_rom[ 1294]='h00000000;
    rd_cycle[ 1295] = 1'b1;  wr_cycle[ 1295] = 1'b0;  addr_rom[ 1295]='h0000003c;  wr_data_rom[ 1295]='h00000000;
    rd_cycle[ 1296] = 1'b1;  wr_cycle[ 1296] = 1'b0;  addr_rom[ 1296]='h00000040;  wr_data_rom[ 1296]='h00000000;
    rd_cycle[ 1297] = 1'b1;  wr_cycle[ 1297] = 1'b0;  addr_rom[ 1297]='h00000044;  wr_data_rom[ 1297]='h00000000;
    rd_cycle[ 1298] = 1'b1;  wr_cycle[ 1298] = 1'b0;  addr_rom[ 1298]='h00000048;  wr_data_rom[ 1298]='h00000000;
    rd_cycle[ 1299] = 1'b1;  wr_cycle[ 1299] = 1'b0;  addr_rom[ 1299]='h0000004c;  wr_data_rom[ 1299]='h00000000;
    rd_cycle[ 1300] = 1'b1;  wr_cycle[ 1300] = 1'b0;  addr_rom[ 1300]='h00000050;  wr_data_rom[ 1300]='h00000000;
    rd_cycle[ 1301] = 1'b1;  wr_cycle[ 1301] = 1'b0;  addr_rom[ 1301]='h00000054;  wr_data_rom[ 1301]='h00000000;
    rd_cycle[ 1302] = 1'b1;  wr_cycle[ 1302] = 1'b0;  addr_rom[ 1302]='h00000058;  wr_data_rom[ 1302]='h00000000;
    rd_cycle[ 1303] = 1'b1;  wr_cycle[ 1303] = 1'b0;  addr_rom[ 1303]='h0000005c;  wr_data_rom[ 1303]='h00000000;
    rd_cycle[ 1304] = 1'b1;  wr_cycle[ 1304] = 1'b0;  addr_rom[ 1304]='h00000060;  wr_data_rom[ 1304]='h00000000;
    rd_cycle[ 1305] = 1'b1;  wr_cycle[ 1305] = 1'b0;  addr_rom[ 1305]='h00000064;  wr_data_rom[ 1305]='h00000000;
    rd_cycle[ 1306] = 1'b1;  wr_cycle[ 1306] = 1'b0;  addr_rom[ 1306]='h00000068;  wr_data_rom[ 1306]='h00000000;
    rd_cycle[ 1307] = 1'b1;  wr_cycle[ 1307] = 1'b0;  addr_rom[ 1307]='h0000006c;  wr_data_rom[ 1307]='h00000000;
    rd_cycle[ 1308] = 1'b1;  wr_cycle[ 1308] = 1'b0;  addr_rom[ 1308]='h00000070;  wr_data_rom[ 1308]='h00000000;
    rd_cycle[ 1309] = 1'b1;  wr_cycle[ 1309] = 1'b0;  addr_rom[ 1309]='h00000074;  wr_data_rom[ 1309]='h00000000;
    rd_cycle[ 1310] = 1'b1;  wr_cycle[ 1310] = 1'b0;  addr_rom[ 1310]='h00000078;  wr_data_rom[ 1310]='h00000000;
    rd_cycle[ 1311] = 1'b1;  wr_cycle[ 1311] = 1'b0;  addr_rom[ 1311]='h0000007c;  wr_data_rom[ 1311]='h00000000;
    rd_cycle[ 1312] = 1'b1;  wr_cycle[ 1312] = 1'b0;  addr_rom[ 1312]='h00000080;  wr_data_rom[ 1312]='h00000000;
    rd_cycle[ 1313] = 1'b1;  wr_cycle[ 1313] = 1'b0;  addr_rom[ 1313]='h00000084;  wr_data_rom[ 1313]='h00000000;
    rd_cycle[ 1314] = 1'b1;  wr_cycle[ 1314] = 1'b0;  addr_rom[ 1314]='h00000088;  wr_data_rom[ 1314]='h00000000;
    rd_cycle[ 1315] = 1'b1;  wr_cycle[ 1315] = 1'b0;  addr_rom[ 1315]='h0000008c;  wr_data_rom[ 1315]='h00000000;
    rd_cycle[ 1316] = 1'b1;  wr_cycle[ 1316] = 1'b0;  addr_rom[ 1316]='h00000090;  wr_data_rom[ 1316]='h00000000;
    rd_cycle[ 1317] = 1'b1;  wr_cycle[ 1317] = 1'b0;  addr_rom[ 1317]='h00000094;  wr_data_rom[ 1317]='h00000000;
    rd_cycle[ 1318] = 1'b1;  wr_cycle[ 1318] = 1'b0;  addr_rom[ 1318]='h00000098;  wr_data_rom[ 1318]='h00000000;
    rd_cycle[ 1319] = 1'b1;  wr_cycle[ 1319] = 1'b0;  addr_rom[ 1319]='h0000009c;  wr_data_rom[ 1319]='h00000000;
    rd_cycle[ 1320] = 1'b1;  wr_cycle[ 1320] = 1'b0;  addr_rom[ 1320]='h000000a0;  wr_data_rom[ 1320]='h00000000;
    rd_cycle[ 1321] = 1'b1;  wr_cycle[ 1321] = 1'b0;  addr_rom[ 1321]='h000000a4;  wr_data_rom[ 1321]='h00000000;
    rd_cycle[ 1322] = 1'b1;  wr_cycle[ 1322] = 1'b0;  addr_rom[ 1322]='h000000a8;  wr_data_rom[ 1322]='h00000000;
    rd_cycle[ 1323] = 1'b1;  wr_cycle[ 1323] = 1'b0;  addr_rom[ 1323]='h000000ac;  wr_data_rom[ 1323]='h00000000;
    rd_cycle[ 1324] = 1'b1;  wr_cycle[ 1324] = 1'b0;  addr_rom[ 1324]='h000000b0;  wr_data_rom[ 1324]='h00000000;
    rd_cycle[ 1325] = 1'b1;  wr_cycle[ 1325] = 1'b0;  addr_rom[ 1325]='h000000b4;  wr_data_rom[ 1325]='h00000000;
    rd_cycle[ 1326] = 1'b1;  wr_cycle[ 1326] = 1'b0;  addr_rom[ 1326]='h000000b8;  wr_data_rom[ 1326]='h00000000;
    rd_cycle[ 1327] = 1'b1;  wr_cycle[ 1327] = 1'b0;  addr_rom[ 1327]='h000000bc;  wr_data_rom[ 1327]='h00000000;
    rd_cycle[ 1328] = 1'b1;  wr_cycle[ 1328] = 1'b0;  addr_rom[ 1328]='h000000c0;  wr_data_rom[ 1328]='h00000000;
    rd_cycle[ 1329] = 1'b1;  wr_cycle[ 1329] = 1'b0;  addr_rom[ 1329]='h000000c4;  wr_data_rom[ 1329]='h00000000;
    rd_cycle[ 1330] = 1'b1;  wr_cycle[ 1330] = 1'b0;  addr_rom[ 1330]='h000000c8;  wr_data_rom[ 1330]='h00000000;
    rd_cycle[ 1331] = 1'b1;  wr_cycle[ 1331] = 1'b0;  addr_rom[ 1331]='h000000cc;  wr_data_rom[ 1331]='h00000000;
    rd_cycle[ 1332] = 1'b1;  wr_cycle[ 1332] = 1'b0;  addr_rom[ 1332]='h000000d0;  wr_data_rom[ 1332]='h00000000;
    rd_cycle[ 1333] = 1'b1;  wr_cycle[ 1333] = 1'b0;  addr_rom[ 1333]='h000000d4;  wr_data_rom[ 1333]='h00000000;
    rd_cycle[ 1334] = 1'b1;  wr_cycle[ 1334] = 1'b0;  addr_rom[ 1334]='h000000d8;  wr_data_rom[ 1334]='h00000000;
    rd_cycle[ 1335] = 1'b1;  wr_cycle[ 1335] = 1'b0;  addr_rom[ 1335]='h000000dc;  wr_data_rom[ 1335]='h00000000;
    rd_cycle[ 1336] = 1'b1;  wr_cycle[ 1336] = 1'b0;  addr_rom[ 1336]='h000000e0;  wr_data_rom[ 1336]='h00000000;
    rd_cycle[ 1337] = 1'b1;  wr_cycle[ 1337] = 1'b0;  addr_rom[ 1337]='h000000e4;  wr_data_rom[ 1337]='h00000000;
    rd_cycle[ 1338] = 1'b1;  wr_cycle[ 1338] = 1'b0;  addr_rom[ 1338]='h000000e8;  wr_data_rom[ 1338]='h00000000;
    rd_cycle[ 1339] = 1'b1;  wr_cycle[ 1339] = 1'b0;  addr_rom[ 1339]='h000000ec;  wr_data_rom[ 1339]='h00000000;
    rd_cycle[ 1340] = 1'b1;  wr_cycle[ 1340] = 1'b0;  addr_rom[ 1340]='h000000f0;  wr_data_rom[ 1340]='h00000000;
    rd_cycle[ 1341] = 1'b1;  wr_cycle[ 1341] = 1'b0;  addr_rom[ 1341]='h000000f4;  wr_data_rom[ 1341]='h00000000;
    rd_cycle[ 1342] = 1'b1;  wr_cycle[ 1342] = 1'b0;  addr_rom[ 1342]='h000000f8;  wr_data_rom[ 1342]='h00000000;
    rd_cycle[ 1343] = 1'b1;  wr_cycle[ 1343] = 1'b0;  addr_rom[ 1343]='h000000fc;  wr_data_rom[ 1343]='h00000000;
    rd_cycle[ 1344] = 1'b1;  wr_cycle[ 1344] = 1'b0;  addr_rom[ 1344]='h00000100;  wr_data_rom[ 1344]='h00000000;
    rd_cycle[ 1345] = 1'b1;  wr_cycle[ 1345] = 1'b0;  addr_rom[ 1345]='h00000104;  wr_data_rom[ 1345]='h00000000;
    rd_cycle[ 1346] = 1'b1;  wr_cycle[ 1346] = 1'b0;  addr_rom[ 1346]='h00000108;  wr_data_rom[ 1346]='h00000000;
    rd_cycle[ 1347] = 1'b1;  wr_cycle[ 1347] = 1'b0;  addr_rom[ 1347]='h0000010c;  wr_data_rom[ 1347]='h00000000;
    rd_cycle[ 1348] = 1'b1;  wr_cycle[ 1348] = 1'b0;  addr_rom[ 1348]='h00000110;  wr_data_rom[ 1348]='h00000000;
    rd_cycle[ 1349] = 1'b1;  wr_cycle[ 1349] = 1'b0;  addr_rom[ 1349]='h00000114;  wr_data_rom[ 1349]='h00000000;
    rd_cycle[ 1350] = 1'b1;  wr_cycle[ 1350] = 1'b0;  addr_rom[ 1350]='h00000118;  wr_data_rom[ 1350]='h00000000;
    rd_cycle[ 1351] = 1'b1;  wr_cycle[ 1351] = 1'b0;  addr_rom[ 1351]='h0000011c;  wr_data_rom[ 1351]='h00000000;
    rd_cycle[ 1352] = 1'b1;  wr_cycle[ 1352] = 1'b0;  addr_rom[ 1352]='h00000120;  wr_data_rom[ 1352]='h00000000;
    rd_cycle[ 1353] = 1'b1;  wr_cycle[ 1353] = 1'b0;  addr_rom[ 1353]='h00000124;  wr_data_rom[ 1353]='h00000000;
    rd_cycle[ 1354] = 1'b1;  wr_cycle[ 1354] = 1'b0;  addr_rom[ 1354]='h00000128;  wr_data_rom[ 1354]='h00000000;
    rd_cycle[ 1355] = 1'b1;  wr_cycle[ 1355] = 1'b0;  addr_rom[ 1355]='h0000012c;  wr_data_rom[ 1355]='h00000000;
    rd_cycle[ 1356] = 1'b1;  wr_cycle[ 1356] = 1'b0;  addr_rom[ 1356]='h00000130;  wr_data_rom[ 1356]='h00000000;
    rd_cycle[ 1357] = 1'b1;  wr_cycle[ 1357] = 1'b0;  addr_rom[ 1357]='h00000134;  wr_data_rom[ 1357]='h00000000;
    rd_cycle[ 1358] = 1'b1;  wr_cycle[ 1358] = 1'b0;  addr_rom[ 1358]='h00000138;  wr_data_rom[ 1358]='h00000000;
    rd_cycle[ 1359] = 1'b1;  wr_cycle[ 1359] = 1'b0;  addr_rom[ 1359]='h0000013c;  wr_data_rom[ 1359]='h00000000;
    rd_cycle[ 1360] = 1'b1;  wr_cycle[ 1360] = 1'b0;  addr_rom[ 1360]='h00000140;  wr_data_rom[ 1360]='h00000000;
    rd_cycle[ 1361] = 1'b1;  wr_cycle[ 1361] = 1'b0;  addr_rom[ 1361]='h00000144;  wr_data_rom[ 1361]='h00000000;
    rd_cycle[ 1362] = 1'b1;  wr_cycle[ 1362] = 1'b0;  addr_rom[ 1362]='h00000148;  wr_data_rom[ 1362]='h00000000;
    rd_cycle[ 1363] = 1'b1;  wr_cycle[ 1363] = 1'b0;  addr_rom[ 1363]='h0000014c;  wr_data_rom[ 1363]='h00000000;
    rd_cycle[ 1364] = 1'b1;  wr_cycle[ 1364] = 1'b0;  addr_rom[ 1364]='h00000150;  wr_data_rom[ 1364]='h00000000;
    rd_cycle[ 1365] = 1'b1;  wr_cycle[ 1365] = 1'b0;  addr_rom[ 1365]='h00000154;  wr_data_rom[ 1365]='h00000000;
    rd_cycle[ 1366] = 1'b1;  wr_cycle[ 1366] = 1'b0;  addr_rom[ 1366]='h00000158;  wr_data_rom[ 1366]='h00000000;
    rd_cycle[ 1367] = 1'b1;  wr_cycle[ 1367] = 1'b0;  addr_rom[ 1367]='h0000015c;  wr_data_rom[ 1367]='h00000000;
    rd_cycle[ 1368] = 1'b1;  wr_cycle[ 1368] = 1'b0;  addr_rom[ 1368]='h00000160;  wr_data_rom[ 1368]='h00000000;
    rd_cycle[ 1369] = 1'b1;  wr_cycle[ 1369] = 1'b0;  addr_rom[ 1369]='h00000164;  wr_data_rom[ 1369]='h00000000;
    rd_cycle[ 1370] = 1'b1;  wr_cycle[ 1370] = 1'b0;  addr_rom[ 1370]='h00000168;  wr_data_rom[ 1370]='h00000000;
    rd_cycle[ 1371] = 1'b1;  wr_cycle[ 1371] = 1'b0;  addr_rom[ 1371]='h0000016c;  wr_data_rom[ 1371]='h00000000;
    rd_cycle[ 1372] = 1'b1;  wr_cycle[ 1372] = 1'b0;  addr_rom[ 1372]='h00000170;  wr_data_rom[ 1372]='h00000000;
    rd_cycle[ 1373] = 1'b1;  wr_cycle[ 1373] = 1'b0;  addr_rom[ 1373]='h00000174;  wr_data_rom[ 1373]='h00000000;
    rd_cycle[ 1374] = 1'b1;  wr_cycle[ 1374] = 1'b0;  addr_rom[ 1374]='h00000178;  wr_data_rom[ 1374]='h00000000;
    rd_cycle[ 1375] = 1'b1;  wr_cycle[ 1375] = 1'b0;  addr_rom[ 1375]='h0000017c;  wr_data_rom[ 1375]='h00000000;
    rd_cycle[ 1376] = 1'b1;  wr_cycle[ 1376] = 1'b0;  addr_rom[ 1376]='h00000180;  wr_data_rom[ 1376]='h00000000;
    rd_cycle[ 1377] = 1'b1;  wr_cycle[ 1377] = 1'b0;  addr_rom[ 1377]='h00000184;  wr_data_rom[ 1377]='h00000000;
    rd_cycle[ 1378] = 1'b1;  wr_cycle[ 1378] = 1'b0;  addr_rom[ 1378]='h00000188;  wr_data_rom[ 1378]='h00000000;
    rd_cycle[ 1379] = 1'b1;  wr_cycle[ 1379] = 1'b0;  addr_rom[ 1379]='h0000018c;  wr_data_rom[ 1379]='h00000000;
    rd_cycle[ 1380] = 1'b1;  wr_cycle[ 1380] = 1'b0;  addr_rom[ 1380]='h00000190;  wr_data_rom[ 1380]='h00000000;
    rd_cycle[ 1381] = 1'b1;  wr_cycle[ 1381] = 1'b0;  addr_rom[ 1381]='h00000194;  wr_data_rom[ 1381]='h00000000;
    rd_cycle[ 1382] = 1'b1;  wr_cycle[ 1382] = 1'b0;  addr_rom[ 1382]='h00000198;  wr_data_rom[ 1382]='h00000000;
    rd_cycle[ 1383] = 1'b1;  wr_cycle[ 1383] = 1'b0;  addr_rom[ 1383]='h0000019c;  wr_data_rom[ 1383]='h00000000;
    rd_cycle[ 1384] = 1'b1;  wr_cycle[ 1384] = 1'b0;  addr_rom[ 1384]='h000001a0;  wr_data_rom[ 1384]='h00000000;
    rd_cycle[ 1385] = 1'b1;  wr_cycle[ 1385] = 1'b0;  addr_rom[ 1385]='h000001a4;  wr_data_rom[ 1385]='h00000000;
    rd_cycle[ 1386] = 1'b1;  wr_cycle[ 1386] = 1'b0;  addr_rom[ 1386]='h000001a8;  wr_data_rom[ 1386]='h00000000;
    rd_cycle[ 1387] = 1'b1;  wr_cycle[ 1387] = 1'b0;  addr_rom[ 1387]='h000001ac;  wr_data_rom[ 1387]='h00000000;
    rd_cycle[ 1388] = 1'b1;  wr_cycle[ 1388] = 1'b0;  addr_rom[ 1388]='h000001b0;  wr_data_rom[ 1388]='h00000000;
    rd_cycle[ 1389] = 1'b1;  wr_cycle[ 1389] = 1'b0;  addr_rom[ 1389]='h000001b4;  wr_data_rom[ 1389]='h00000000;
    rd_cycle[ 1390] = 1'b1;  wr_cycle[ 1390] = 1'b0;  addr_rom[ 1390]='h000001b8;  wr_data_rom[ 1390]='h00000000;
    rd_cycle[ 1391] = 1'b1;  wr_cycle[ 1391] = 1'b0;  addr_rom[ 1391]='h000001bc;  wr_data_rom[ 1391]='h00000000;
    rd_cycle[ 1392] = 1'b1;  wr_cycle[ 1392] = 1'b0;  addr_rom[ 1392]='h000001c0;  wr_data_rom[ 1392]='h00000000;
    rd_cycle[ 1393] = 1'b1;  wr_cycle[ 1393] = 1'b0;  addr_rom[ 1393]='h000001c4;  wr_data_rom[ 1393]='h00000000;
    rd_cycle[ 1394] = 1'b1;  wr_cycle[ 1394] = 1'b0;  addr_rom[ 1394]='h000001c8;  wr_data_rom[ 1394]='h00000000;
    rd_cycle[ 1395] = 1'b1;  wr_cycle[ 1395] = 1'b0;  addr_rom[ 1395]='h000001cc;  wr_data_rom[ 1395]='h00000000;
    rd_cycle[ 1396] = 1'b1;  wr_cycle[ 1396] = 1'b0;  addr_rom[ 1396]='h000001d0;  wr_data_rom[ 1396]='h00000000;
    rd_cycle[ 1397] = 1'b1;  wr_cycle[ 1397] = 1'b0;  addr_rom[ 1397]='h000001d4;  wr_data_rom[ 1397]='h00000000;
    rd_cycle[ 1398] = 1'b1;  wr_cycle[ 1398] = 1'b0;  addr_rom[ 1398]='h000001d8;  wr_data_rom[ 1398]='h00000000;
    rd_cycle[ 1399] = 1'b1;  wr_cycle[ 1399] = 1'b0;  addr_rom[ 1399]='h000001dc;  wr_data_rom[ 1399]='h00000000;
    rd_cycle[ 1400] = 1'b1;  wr_cycle[ 1400] = 1'b0;  addr_rom[ 1400]='h000001e0;  wr_data_rom[ 1400]='h00000000;
    rd_cycle[ 1401] = 1'b1;  wr_cycle[ 1401] = 1'b0;  addr_rom[ 1401]='h000001e4;  wr_data_rom[ 1401]='h00000000;
    rd_cycle[ 1402] = 1'b1;  wr_cycle[ 1402] = 1'b0;  addr_rom[ 1402]='h000001e8;  wr_data_rom[ 1402]='h00000000;
    rd_cycle[ 1403] = 1'b1;  wr_cycle[ 1403] = 1'b0;  addr_rom[ 1403]='h000001ec;  wr_data_rom[ 1403]='h00000000;
    rd_cycle[ 1404] = 1'b1;  wr_cycle[ 1404] = 1'b0;  addr_rom[ 1404]='h000001f0;  wr_data_rom[ 1404]='h00000000;
    rd_cycle[ 1405] = 1'b1;  wr_cycle[ 1405] = 1'b0;  addr_rom[ 1405]='h000001f4;  wr_data_rom[ 1405]='h00000000;
    rd_cycle[ 1406] = 1'b1;  wr_cycle[ 1406] = 1'b0;  addr_rom[ 1406]='h000001f8;  wr_data_rom[ 1406]='h00000000;
    rd_cycle[ 1407] = 1'b1;  wr_cycle[ 1407] = 1'b0;  addr_rom[ 1407]='h000001fc;  wr_data_rom[ 1407]='h00000000;
    rd_cycle[ 1408] = 1'b1;  wr_cycle[ 1408] = 1'b0;  addr_rom[ 1408]='h00000200;  wr_data_rom[ 1408]='h00000000;
    rd_cycle[ 1409] = 1'b1;  wr_cycle[ 1409] = 1'b0;  addr_rom[ 1409]='h00000204;  wr_data_rom[ 1409]='h00000000;
    rd_cycle[ 1410] = 1'b1;  wr_cycle[ 1410] = 1'b0;  addr_rom[ 1410]='h00000208;  wr_data_rom[ 1410]='h00000000;
    rd_cycle[ 1411] = 1'b1;  wr_cycle[ 1411] = 1'b0;  addr_rom[ 1411]='h0000020c;  wr_data_rom[ 1411]='h00000000;
    rd_cycle[ 1412] = 1'b1;  wr_cycle[ 1412] = 1'b0;  addr_rom[ 1412]='h00000210;  wr_data_rom[ 1412]='h00000000;
    rd_cycle[ 1413] = 1'b1;  wr_cycle[ 1413] = 1'b0;  addr_rom[ 1413]='h00000214;  wr_data_rom[ 1413]='h00000000;
    rd_cycle[ 1414] = 1'b1;  wr_cycle[ 1414] = 1'b0;  addr_rom[ 1414]='h00000218;  wr_data_rom[ 1414]='h00000000;
    rd_cycle[ 1415] = 1'b1;  wr_cycle[ 1415] = 1'b0;  addr_rom[ 1415]='h0000021c;  wr_data_rom[ 1415]='h00000000;
    rd_cycle[ 1416] = 1'b1;  wr_cycle[ 1416] = 1'b0;  addr_rom[ 1416]='h00000220;  wr_data_rom[ 1416]='h00000000;
    rd_cycle[ 1417] = 1'b1;  wr_cycle[ 1417] = 1'b0;  addr_rom[ 1417]='h00000224;  wr_data_rom[ 1417]='h00000000;
    rd_cycle[ 1418] = 1'b1;  wr_cycle[ 1418] = 1'b0;  addr_rom[ 1418]='h00000228;  wr_data_rom[ 1418]='h00000000;
    rd_cycle[ 1419] = 1'b1;  wr_cycle[ 1419] = 1'b0;  addr_rom[ 1419]='h0000022c;  wr_data_rom[ 1419]='h00000000;
    rd_cycle[ 1420] = 1'b1;  wr_cycle[ 1420] = 1'b0;  addr_rom[ 1420]='h00000230;  wr_data_rom[ 1420]='h00000000;
    rd_cycle[ 1421] = 1'b1;  wr_cycle[ 1421] = 1'b0;  addr_rom[ 1421]='h00000234;  wr_data_rom[ 1421]='h00000000;
    rd_cycle[ 1422] = 1'b1;  wr_cycle[ 1422] = 1'b0;  addr_rom[ 1422]='h00000238;  wr_data_rom[ 1422]='h00000000;
    rd_cycle[ 1423] = 1'b1;  wr_cycle[ 1423] = 1'b0;  addr_rom[ 1423]='h0000023c;  wr_data_rom[ 1423]='h00000000;
    rd_cycle[ 1424] = 1'b1;  wr_cycle[ 1424] = 1'b0;  addr_rom[ 1424]='h00000240;  wr_data_rom[ 1424]='h00000000;
    rd_cycle[ 1425] = 1'b1;  wr_cycle[ 1425] = 1'b0;  addr_rom[ 1425]='h00000244;  wr_data_rom[ 1425]='h00000000;
    rd_cycle[ 1426] = 1'b1;  wr_cycle[ 1426] = 1'b0;  addr_rom[ 1426]='h00000248;  wr_data_rom[ 1426]='h00000000;
    rd_cycle[ 1427] = 1'b1;  wr_cycle[ 1427] = 1'b0;  addr_rom[ 1427]='h0000024c;  wr_data_rom[ 1427]='h00000000;
    rd_cycle[ 1428] = 1'b1;  wr_cycle[ 1428] = 1'b0;  addr_rom[ 1428]='h00000250;  wr_data_rom[ 1428]='h00000000;
    rd_cycle[ 1429] = 1'b1;  wr_cycle[ 1429] = 1'b0;  addr_rom[ 1429]='h00000254;  wr_data_rom[ 1429]='h00000000;
    rd_cycle[ 1430] = 1'b1;  wr_cycle[ 1430] = 1'b0;  addr_rom[ 1430]='h00000258;  wr_data_rom[ 1430]='h00000000;
    rd_cycle[ 1431] = 1'b1;  wr_cycle[ 1431] = 1'b0;  addr_rom[ 1431]='h0000025c;  wr_data_rom[ 1431]='h00000000;
    rd_cycle[ 1432] = 1'b1;  wr_cycle[ 1432] = 1'b0;  addr_rom[ 1432]='h00000260;  wr_data_rom[ 1432]='h00000000;
    rd_cycle[ 1433] = 1'b1;  wr_cycle[ 1433] = 1'b0;  addr_rom[ 1433]='h00000264;  wr_data_rom[ 1433]='h00000000;
    rd_cycle[ 1434] = 1'b1;  wr_cycle[ 1434] = 1'b0;  addr_rom[ 1434]='h00000268;  wr_data_rom[ 1434]='h00000000;
    rd_cycle[ 1435] = 1'b1;  wr_cycle[ 1435] = 1'b0;  addr_rom[ 1435]='h0000026c;  wr_data_rom[ 1435]='h00000000;
    rd_cycle[ 1436] = 1'b1;  wr_cycle[ 1436] = 1'b0;  addr_rom[ 1436]='h00000270;  wr_data_rom[ 1436]='h00000000;
    rd_cycle[ 1437] = 1'b1;  wr_cycle[ 1437] = 1'b0;  addr_rom[ 1437]='h00000274;  wr_data_rom[ 1437]='h00000000;
    rd_cycle[ 1438] = 1'b1;  wr_cycle[ 1438] = 1'b0;  addr_rom[ 1438]='h00000278;  wr_data_rom[ 1438]='h00000000;
    rd_cycle[ 1439] = 1'b1;  wr_cycle[ 1439] = 1'b0;  addr_rom[ 1439]='h0000027c;  wr_data_rom[ 1439]='h00000000;
    rd_cycle[ 1440] = 1'b1;  wr_cycle[ 1440] = 1'b0;  addr_rom[ 1440]='h00000280;  wr_data_rom[ 1440]='h00000000;
    rd_cycle[ 1441] = 1'b1;  wr_cycle[ 1441] = 1'b0;  addr_rom[ 1441]='h00000284;  wr_data_rom[ 1441]='h00000000;
    rd_cycle[ 1442] = 1'b1;  wr_cycle[ 1442] = 1'b0;  addr_rom[ 1442]='h00000288;  wr_data_rom[ 1442]='h00000000;
    rd_cycle[ 1443] = 1'b1;  wr_cycle[ 1443] = 1'b0;  addr_rom[ 1443]='h0000028c;  wr_data_rom[ 1443]='h00000000;
    rd_cycle[ 1444] = 1'b1;  wr_cycle[ 1444] = 1'b0;  addr_rom[ 1444]='h00000290;  wr_data_rom[ 1444]='h00000000;
    rd_cycle[ 1445] = 1'b1;  wr_cycle[ 1445] = 1'b0;  addr_rom[ 1445]='h00000294;  wr_data_rom[ 1445]='h00000000;
    rd_cycle[ 1446] = 1'b1;  wr_cycle[ 1446] = 1'b0;  addr_rom[ 1446]='h00000298;  wr_data_rom[ 1446]='h00000000;
    rd_cycle[ 1447] = 1'b1;  wr_cycle[ 1447] = 1'b0;  addr_rom[ 1447]='h0000029c;  wr_data_rom[ 1447]='h00000000;
    rd_cycle[ 1448] = 1'b1;  wr_cycle[ 1448] = 1'b0;  addr_rom[ 1448]='h000002a0;  wr_data_rom[ 1448]='h00000000;
    rd_cycle[ 1449] = 1'b1;  wr_cycle[ 1449] = 1'b0;  addr_rom[ 1449]='h000002a4;  wr_data_rom[ 1449]='h00000000;
    rd_cycle[ 1450] = 1'b1;  wr_cycle[ 1450] = 1'b0;  addr_rom[ 1450]='h000002a8;  wr_data_rom[ 1450]='h00000000;
    rd_cycle[ 1451] = 1'b1;  wr_cycle[ 1451] = 1'b0;  addr_rom[ 1451]='h000002ac;  wr_data_rom[ 1451]='h00000000;
    rd_cycle[ 1452] = 1'b1;  wr_cycle[ 1452] = 1'b0;  addr_rom[ 1452]='h000002b0;  wr_data_rom[ 1452]='h00000000;
    rd_cycle[ 1453] = 1'b1;  wr_cycle[ 1453] = 1'b0;  addr_rom[ 1453]='h000002b4;  wr_data_rom[ 1453]='h00000000;
    rd_cycle[ 1454] = 1'b1;  wr_cycle[ 1454] = 1'b0;  addr_rom[ 1454]='h000002b8;  wr_data_rom[ 1454]='h00000000;
    rd_cycle[ 1455] = 1'b1;  wr_cycle[ 1455] = 1'b0;  addr_rom[ 1455]='h000002bc;  wr_data_rom[ 1455]='h00000000;
    rd_cycle[ 1456] = 1'b1;  wr_cycle[ 1456] = 1'b0;  addr_rom[ 1456]='h000002c0;  wr_data_rom[ 1456]='h00000000;
    rd_cycle[ 1457] = 1'b1;  wr_cycle[ 1457] = 1'b0;  addr_rom[ 1457]='h000002c4;  wr_data_rom[ 1457]='h00000000;
    rd_cycle[ 1458] = 1'b1;  wr_cycle[ 1458] = 1'b0;  addr_rom[ 1458]='h000002c8;  wr_data_rom[ 1458]='h00000000;
    rd_cycle[ 1459] = 1'b1;  wr_cycle[ 1459] = 1'b0;  addr_rom[ 1459]='h000002cc;  wr_data_rom[ 1459]='h00000000;
    rd_cycle[ 1460] = 1'b1;  wr_cycle[ 1460] = 1'b0;  addr_rom[ 1460]='h000002d0;  wr_data_rom[ 1460]='h00000000;
    rd_cycle[ 1461] = 1'b1;  wr_cycle[ 1461] = 1'b0;  addr_rom[ 1461]='h000002d4;  wr_data_rom[ 1461]='h00000000;
    rd_cycle[ 1462] = 1'b1;  wr_cycle[ 1462] = 1'b0;  addr_rom[ 1462]='h000002d8;  wr_data_rom[ 1462]='h00000000;
    rd_cycle[ 1463] = 1'b1;  wr_cycle[ 1463] = 1'b0;  addr_rom[ 1463]='h000002dc;  wr_data_rom[ 1463]='h00000000;
    rd_cycle[ 1464] = 1'b1;  wr_cycle[ 1464] = 1'b0;  addr_rom[ 1464]='h000002e0;  wr_data_rom[ 1464]='h00000000;
    rd_cycle[ 1465] = 1'b1;  wr_cycle[ 1465] = 1'b0;  addr_rom[ 1465]='h000002e4;  wr_data_rom[ 1465]='h00000000;
    rd_cycle[ 1466] = 1'b1;  wr_cycle[ 1466] = 1'b0;  addr_rom[ 1466]='h000002e8;  wr_data_rom[ 1466]='h00000000;
    rd_cycle[ 1467] = 1'b1;  wr_cycle[ 1467] = 1'b0;  addr_rom[ 1467]='h000002ec;  wr_data_rom[ 1467]='h00000000;
    rd_cycle[ 1468] = 1'b1;  wr_cycle[ 1468] = 1'b0;  addr_rom[ 1468]='h000002f0;  wr_data_rom[ 1468]='h00000000;
    rd_cycle[ 1469] = 1'b1;  wr_cycle[ 1469] = 1'b0;  addr_rom[ 1469]='h000002f4;  wr_data_rom[ 1469]='h00000000;
    rd_cycle[ 1470] = 1'b1;  wr_cycle[ 1470] = 1'b0;  addr_rom[ 1470]='h000002f8;  wr_data_rom[ 1470]='h00000000;
    rd_cycle[ 1471] = 1'b1;  wr_cycle[ 1471] = 1'b0;  addr_rom[ 1471]='h000002fc;  wr_data_rom[ 1471]='h00000000;
    rd_cycle[ 1472] = 1'b1;  wr_cycle[ 1472] = 1'b0;  addr_rom[ 1472]='h00000300;  wr_data_rom[ 1472]='h00000000;
    rd_cycle[ 1473] = 1'b1;  wr_cycle[ 1473] = 1'b0;  addr_rom[ 1473]='h00000304;  wr_data_rom[ 1473]='h00000000;
    rd_cycle[ 1474] = 1'b1;  wr_cycle[ 1474] = 1'b0;  addr_rom[ 1474]='h00000308;  wr_data_rom[ 1474]='h00000000;
    rd_cycle[ 1475] = 1'b1;  wr_cycle[ 1475] = 1'b0;  addr_rom[ 1475]='h0000030c;  wr_data_rom[ 1475]='h00000000;
    rd_cycle[ 1476] = 1'b1;  wr_cycle[ 1476] = 1'b0;  addr_rom[ 1476]='h00000310;  wr_data_rom[ 1476]='h00000000;
    rd_cycle[ 1477] = 1'b1;  wr_cycle[ 1477] = 1'b0;  addr_rom[ 1477]='h00000314;  wr_data_rom[ 1477]='h00000000;
    rd_cycle[ 1478] = 1'b1;  wr_cycle[ 1478] = 1'b0;  addr_rom[ 1478]='h00000318;  wr_data_rom[ 1478]='h00000000;
    rd_cycle[ 1479] = 1'b1;  wr_cycle[ 1479] = 1'b0;  addr_rom[ 1479]='h0000031c;  wr_data_rom[ 1479]='h00000000;
    rd_cycle[ 1480] = 1'b1;  wr_cycle[ 1480] = 1'b0;  addr_rom[ 1480]='h00000320;  wr_data_rom[ 1480]='h00000000;
    rd_cycle[ 1481] = 1'b1;  wr_cycle[ 1481] = 1'b0;  addr_rom[ 1481]='h00000324;  wr_data_rom[ 1481]='h00000000;
    rd_cycle[ 1482] = 1'b1;  wr_cycle[ 1482] = 1'b0;  addr_rom[ 1482]='h00000328;  wr_data_rom[ 1482]='h00000000;
    rd_cycle[ 1483] = 1'b1;  wr_cycle[ 1483] = 1'b0;  addr_rom[ 1483]='h0000032c;  wr_data_rom[ 1483]='h00000000;
    rd_cycle[ 1484] = 1'b1;  wr_cycle[ 1484] = 1'b0;  addr_rom[ 1484]='h00000330;  wr_data_rom[ 1484]='h00000000;
    rd_cycle[ 1485] = 1'b1;  wr_cycle[ 1485] = 1'b0;  addr_rom[ 1485]='h00000334;  wr_data_rom[ 1485]='h00000000;
    rd_cycle[ 1486] = 1'b1;  wr_cycle[ 1486] = 1'b0;  addr_rom[ 1486]='h00000338;  wr_data_rom[ 1486]='h00000000;
    rd_cycle[ 1487] = 1'b1;  wr_cycle[ 1487] = 1'b0;  addr_rom[ 1487]='h0000033c;  wr_data_rom[ 1487]='h00000000;
    rd_cycle[ 1488] = 1'b1;  wr_cycle[ 1488] = 1'b0;  addr_rom[ 1488]='h00000340;  wr_data_rom[ 1488]='h00000000;
    rd_cycle[ 1489] = 1'b1;  wr_cycle[ 1489] = 1'b0;  addr_rom[ 1489]='h00000344;  wr_data_rom[ 1489]='h00000000;
    rd_cycle[ 1490] = 1'b1;  wr_cycle[ 1490] = 1'b0;  addr_rom[ 1490]='h00000348;  wr_data_rom[ 1490]='h00000000;
    rd_cycle[ 1491] = 1'b1;  wr_cycle[ 1491] = 1'b0;  addr_rom[ 1491]='h0000034c;  wr_data_rom[ 1491]='h00000000;
    rd_cycle[ 1492] = 1'b1;  wr_cycle[ 1492] = 1'b0;  addr_rom[ 1492]='h00000350;  wr_data_rom[ 1492]='h00000000;
    rd_cycle[ 1493] = 1'b1;  wr_cycle[ 1493] = 1'b0;  addr_rom[ 1493]='h00000354;  wr_data_rom[ 1493]='h00000000;
    rd_cycle[ 1494] = 1'b1;  wr_cycle[ 1494] = 1'b0;  addr_rom[ 1494]='h00000358;  wr_data_rom[ 1494]='h00000000;
    rd_cycle[ 1495] = 1'b1;  wr_cycle[ 1495] = 1'b0;  addr_rom[ 1495]='h0000035c;  wr_data_rom[ 1495]='h00000000;
    rd_cycle[ 1496] = 1'b1;  wr_cycle[ 1496] = 1'b0;  addr_rom[ 1496]='h00000360;  wr_data_rom[ 1496]='h00000000;
    rd_cycle[ 1497] = 1'b1;  wr_cycle[ 1497] = 1'b0;  addr_rom[ 1497]='h00000364;  wr_data_rom[ 1497]='h00000000;
    rd_cycle[ 1498] = 1'b1;  wr_cycle[ 1498] = 1'b0;  addr_rom[ 1498]='h00000368;  wr_data_rom[ 1498]='h00000000;
    rd_cycle[ 1499] = 1'b1;  wr_cycle[ 1499] = 1'b0;  addr_rom[ 1499]='h0000036c;  wr_data_rom[ 1499]='h00000000;
    rd_cycle[ 1500] = 1'b1;  wr_cycle[ 1500] = 1'b0;  addr_rom[ 1500]='h00000370;  wr_data_rom[ 1500]='h00000000;
    rd_cycle[ 1501] = 1'b1;  wr_cycle[ 1501] = 1'b0;  addr_rom[ 1501]='h00000374;  wr_data_rom[ 1501]='h00000000;
    rd_cycle[ 1502] = 1'b1;  wr_cycle[ 1502] = 1'b0;  addr_rom[ 1502]='h00000378;  wr_data_rom[ 1502]='h00000000;
    rd_cycle[ 1503] = 1'b1;  wr_cycle[ 1503] = 1'b0;  addr_rom[ 1503]='h0000037c;  wr_data_rom[ 1503]='h00000000;
    rd_cycle[ 1504] = 1'b1;  wr_cycle[ 1504] = 1'b0;  addr_rom[ 1504]='h00000380;  wr_data_rom[ 1504]='h00000000;
    rd_cycle[ 1505] = 1'b1;  wr_cycle[ 1505] = 1'b0;  addr_rom[ 1505]='h00000384;  wr_data_rom[ 1505]='h00000000;
    rd_cycle[ 1506] = 1'b1;  wr_cycle[ 1506] = 1'b0;  addr_rom[ 1506]='h00000388;  wr_data_rom[ 1506]='h00000000;
    rd_cycle[ 1507] = 1'b1;  wr_cycle[ 1507] = 1'b0;  addr_rom[ 1507]='h0000038c;  wr_data_rom[ 1507]='h00000000;
    rd_cycle[ 1508] = 1'b1;  wr_cycle[ 1508] = 1'b0;  addr_rom[ 1508]='h00000390;  wr_data_rom[ 1508]='h00000000;
    rd_cycle[ 1509] = 1'b1;  wr_cycle[ 1509] = 1'b0;  addr_rom[ 1509]='h00000394;  wr_data_rom[ 1509]='h00000000;
    rd_cycle[ 1510] = 1'b1;  wr_cycle[ 1510] = 1'b0;  addr_rom[ 1510]='h00000398;  wr_data_rom[ 1510]='h00000000;
    rd_cycle[ 1511] = 1'b1;  wr_cycle[ 1511] = 1'b0;  addr_rom[ 1511]='h0000039c;  wr_data_rom[ 1511]='h00000000;
    rd_cycle[ 1512] = 1'b1;  wr_cycle[ 1512] = 1'b0;  addr_rom[ 1512]='h000003a0;  wr_data_rom[ 1512]='h00000000;
    rd_cycle[ 1513] = 1'b1;  wr_cycle[ 1513] = 1'b0;  addr_rom[ 1513]='h000003a4;  wr_data_rom[ 1513]='h00000000;
    rd_cycle[ 1514] = 1'b1;  wr_cycle[ 1514] = 1'b0;  addr_rom[ 1514]='h000003a8;  wr_data_rom[ 1514]='h00000000;
    rd_cycle[ 1515] = 1'b1;  wr_cycle[ 1515] = 1'b0;  addr_rom[ 1515]='h000003ac;  wr_data_rom[ 1515]='h00000000;
    rd_cycle[ 1516] = 1'b1;  wr_cycle[ 1516] = 1'b0;  addr_rom[ 1516]='h000003b0;  wr_data_rom[ 1516]='h00000000;
    rd_cycle[ 1517] = 1'b1;  wr_cycle[ 1517] = 1'b0;  addr_rom[ 1517]='h000003b4;  wr_data_rom[ 1517]='h00000000;
    rd_cycle[ 1518] = 1'b1;  wr_cycle[ 1518] = 1'b0;  addr_rom[ 1518]='h000003b8;  wr_data_rom[ 1518]='h00000000;
    rd_cycle[ 1519] = 1'b1;  wr_cycle[ 1519] = 1'b0;  addr_rom[ 1519]='h000003bc;  wr_data_rom[ 1519]='h00000000;
    rd_cycle[ 1520] = 1'b1;  wr_cycle[ 1520] = 1'b0;  addr_rom[ 1520]='h000003c0;  wr_data_rom[ 1520]='h00000000;
    rd_cycle[ 1521] = 1'b1;  wr_cycle[ 1521] = 1'b0;  addr_rom[ 1521]='h000003c4;  wr_data_rom[ 1521]='h00000000;
    rd_cycle[ 1522] = 1'b1;  wr_cycle[ 1522] = 1'b0;  addr_rom[ 1522]='h000003c8;  wr_data_rom[ 1522]='h00000000;
    rd_cycle[ 1523] = 1'b1;  wr_cycle[ 1523] = 1'b0;  addr_rom[ 1523]='h000003cc;  wr_data_rom[ 1523]='h00000000;
    rd_cycle[ 1524] = 1'b1;  wr_cycle[ 1524] = 1'b0;  addr_rom[ 1524]='h000003d0;  wr_data_rom[ 1524]='h00000000;
    rd_cycle[ 1525] = 1'b1;  wr_cycle[ 1525] = 1'b0;  addr_rom[ 1525]='h000003d4;  wr_data_rom[ 1525]='h00000000;
    rd_cycle[ 1526] = 1'b1;  wr_cycle[ 1526] = 1'b0;  addr_rom[ 1526]='h000003d8;  wr_data_rom[ 1526]='h00000000;
    rd_cycle[ 1527] = 1'b1;  wr_cycle[ 1527] = 1'b0;  addr_rom[ 1527]='h000003dc;  wr_data_rom[ 1527]='h00000000;
    rd_cycle[ 1528] = 1'b1;  wr_cycle[ 1528] = 1'b0;  addr_rom[ 1528]='h000003e0;  wr_data_rom[ 1528]='h00000000;
    rd_cycle[ 1529] = 1'b1;  wr_cycle[ 1529] = 1'b0;  addr_rom[ 1529]='h000003e4;  wr_data_rom[ 1529]='h00000000;
    rd_cycle[ 1530] = 1'b1;  wr_cycle[ 1530] = 1'b0;  addr_rom[ 1530]='h000003e8;  wr_data_rom[ 1530]='h00000000;
    rd_cycle[ 1531] = 1'b1;  wr_cycle[ 1531] = 1'b0;  addr_rom[ 1531]='h000003ec;  wr_data_rom[ 1531]='h00000000;
    rd_cycle[ 1532] = 1'b1;  wr_cycle[ 1532] = 1'b0;  addr_rom[ 1532]='h000003f0;  wr_data_rom[ 1532]='h00000000;
    rd_cycle[ 1533] = 1'b1;  wr_cycle[ 1533] = 1'b0;  addr_rom[ 1533]='h000003f4;  wr_data_rom[ 1533]='h00000000;
    rd_cycle[ 1534] = 1'b1;  wr_cycle[ 1534] = 1'b0;  addr_rom[ 1534]='h000003f8;  wr_data_rom[ 1534]='h00000000;
    rd_cycle[ 1535] = 1'b1;  wr_cycle[ 1535] = 1'b0;  addr_rom[ 1535]='h000003fc;  wr_data_rom[ 1535]='h00000000;
end

initial begin
    validation_data[    0] = 'h000001a9; 
    validation_data[    1] = 'h000003c0; 
    validation_data[    2] = 'h00000237; 
    validation_data[    3] = 'h0000018b; 
    validation_data[    4] = 'h0000034f; 
    validation_data[    5] = 'h000001bf; 
    validation_data[    6] = 'h00000262; 
    validation_data[    7] = 'h0000036a; 
    validation_data[    8] = 'h00000157; 
    validation_data[    9] = 'h0000005f; 
    validation_data[   10] = 'h000002de; 
    validation_data[   11] = 'h00000325; 
    validation_data[   12] = 'h000000ac; 
    validation_data[   13] = 'h00000308; 
    validation_data[   14] = 'h000002bf; 
    validation_data[   15] = 'h00000332; 
    validation_data[   16] = 'h000001d2; 
    validation_data[   17] = 'h000002b1; 
    validation_data[   18] = 'h00000231; 
    validation_data[   19] = 'h000000ca; 
    validation_data[   20] = 'h00000041; 
    validation_data[   21] = 'h0000011c; 
    validation_data[   22] = 'h000003e7; 
    validation_data[   23] = 'h0000033e; 
    validation_data[   24] = 'h00000388; 
    validation_data[   25] = 'h00000042; 
    validation_data[   26] = 'h000000c4; 
    validation_data[   27] = 'h000001a3; 
    validation_data[   28] = 'h00000189; 
    validation_data[   29] = 'h000001b9; 
    validation_data[   30] = 'h00000028; 
    validation_data[   31] = 'h000000eb; 
    validation_data[   32] = 'h000000af; 
    validation_data[   33] = 'h00000286; 
    validation_data[   34] = 'h000000ca; 
    validation_data[   35] = 'h00000142; 
    validation_data[   36] = 'h00000220; 
    validation_data[   37] = 'h000002b9; 
    validation_data[   38] = 'h00000014; 
    validation_data[   39] = 'h000002c1; 
    validation_data[   40] = 'h0000013c; 
    validation_data[   41] = 'h00000321; 
    validation_data[   42] = 'h00000130; 
    validation_data[   43] = 'h00000144; 
    validation_data[   44] = 'h00000305; 
    validation_data[   45] = 'h0000025e; 
    validation_data[   46] = 'h000002f6; 
    validation_data[   47] = 'h000001d7; 
    validation_data[   48] = 'h000001b4; 
    validation_data[   49] = 'h0000015e; 
    validation_data[   50] = 'h0000001c; 
    validation_data[   51] = 'h000000b8; 
    validation_data[   52] = 'h000001f5; 
    validation_data[   53] = 'h000003f7; 
    validation_data[   54] = 'h000002fc; 
    validation_data[   55] = 'h000003f1; 
    validation_data[   56] = 'h00000361; 
    validation_data[   57] = 'h000003d4; 
    validation_data[   58] = 'h0000009b; 
    validation_data[   59] = 'h00000293; 
    validation_data[   60] = 'h00000261; 
    validation_data[   61] = 'h0000036f; 
    validation_data[   62] = 'h000002c2; 
    validation_data[   63] = 'h00000171; 
    validation_data[   64] = 'h00000176; 
    validation_data[   65] = 'h000001a2; 
    validation_data[   66] = 'h0000003e; 
    validation_data[   67] = 'h00000209; 
    validation_data[   68] = 'h00000259; 
    validation_data[   69] = 'h00000384; 
    validation_data[   70] = 'h000003e0; 
    validation_data[   71] = 'h00000338; 
    validation_data[   72] = 'h00000314; 
    validation_data[   73] = 'h000001b8; 
    validation_data[   74] = 'h00000325; 
    validation_data[   75] = 'h00000163; 
    validation_data[   76] = 'h0000000e; 
    validation_data[   77] = 'h000001ed; 
    validation_data[   78] = 'h000000db; 
    validation_data[   79] = 'h00000224; 
    validation_data[   80] = 'h000000bd; 
    validation_data[   81] = 'h00000327; 
    validation_data[   82] = 'h00000367; 
    validation_data[   83] = 'h00000130; 
    validation_data[   84] = 'h000003ed; 
    validation_data[   85] = 'h00000233; 
    validation_data[   86] = 'h0000036c; 
    validation_data[   87] = 'h000003f8; 
    validation_data[   88] = 'h0000033a; 
    validation_data[   89] = 'h000001eb; 
    validation_data[   90] = 'h00000052; 
    validation_data[   91] = 'h000000ea; 
    validation_data[   92] = 'h0000027f; 
    validation_data[   93] = 'h000002b0; 
    validation_data[   94] = 'h0000012f; 
    validation_data[   95] = 'h00000107; 
    validation_data[   96] = 'h000003c2; 
    validation_data[   97] = 'h0000003c; 
    validation_data[   98] = 'h00000053; 
    validation_data[   99] = 'h0000034b; 
    validation_data[  100] = 'h00000059; 
    validation_data[  101] = 'h00000318; 
    validation_data[  102] = 'h000001f8; 
    validation_data[  103] = 'h000003d5; 
    validation_data[  104] = 'h000000b5; 
    validation_data[  105] = 'h0000026a; 
    validation_data[  106] = 'h000002f5; 
    validation_data[  107] = 'h0000000a; 
    validation_data[  108] = 'h000003fd; 
    validation_data[  109] = 'h00000350; 
    validation_data[  110] = 'h00000304; 
    validation_data[  111] = 'h00000070; 
    validation_data[  112] = 'h00000379; 
    validation_data[  113] = 'h000003d4; 
    validation_data[  114] = 'h00000366; 
    validation_data[  115] = 'h00000189; 
    validation_data[  116] = 'h00000040; 
    validation_data[  117] = 'h00000028; 
    validation_data[  118] = 'h00000130; 
    validation_data[  119] = 'h000002e0; 
    validation_data[  120] = 'h00000105; 
    validation_data[  121] = 'h000000d0; 
    validation_data[  122] = 'h00000058; 
    validation_data[  123] = 'h0000034e; 
    validation_data[  124] = 'h00000154; 
    validation_data[  125] = 'h00000279; 
    validation_data[  126] = 'h0000018b; 
    validation_data[  127] = 'h00000182; 
    validation_data[  128] = 'h00000317; 
    validation_data[  129] = 'h00000365; 
    validation_data[  130] = 'h000000f1; 
    validation_data[  131] = 'h0000010b; 
    validation_data[  132] = 'h000000a5; 
    validation_data[  133] = 'h00000331; 
    validation_data[  134] = 'h00000266; 
    validation_data[  135] = 'h000003f9; 
    validation_data[  136] = 'h000000ca; 
    validation_data[  137] = 'h000000bb; 
    validation_data[  138] = 'h0000017d; 
    validation_data[  139] = 'h00000141; 
    validation_data[  140] = 'h00000371; 
    validation_data[  141] = 'h000000d9; 
    validation_data[  142] = 'h000003f0; 
    validation_data[  143] = 'h00000328; 
    validation_data[  144] = 'h000001e6; 
    validation_data[  145] = 'h00000159; 
    validation_data[  146] = 'h000000a4; 
    validation_data[  147] = 'h000001c5; 
    validation_data[  148] = 'h00000125; 
    validation_data[  149] = 'h000001a1; 
    validation_data[  150] = 'h000001a1; 
    validation_data[  151] = 'h00000311; 
    validation_data[  152] = 'h000000dd; 
    validation_data[  153] = 'h000002f7; 
    validation_data[  154] = 'h0000001f; 
    validation_data[  155] = 'h0000038b; 
    validation_data[  156] = 'h0000028b; 
    validation_data[  157] = 'h000002dc; 
    validation_data[  158] = 'h00000094; 
    validation_data[  159] = 'h00000101; 
    validation_data[  160] = 'h00000074; 
    validation_data[  161] = 'h000000dd; 
    validation_data[  162] = 'h000003ef; 
    validation_data[  163] = 'h000003af; 
    validation_data[  164] = 'h000003fc; 
    validation_data[  165] = 'h00000354; 
    validation_data[  166] = 'h000000e4; 
    validation_data[  167] = 'h00000140; 
    validation_data[  168] = 'h0000008e; 
    validation_data[  169] = 'h00000106; 
    validation_data[  170] = 'h00000011; 
    validation_data[  171] = 'h000001f1; 
    validation_data[  172] = 'h0000036a; 
    validation_data[  173] = 'h00000004; 
    validation_data[  174] = 'h000002e0; 
    validation_data[  175] = 'h0000003a; 
    validation_data[  176] = 'h00000224; 
    validation_data[  177] = 'h000001dc; 
    validation_data[  178] = 'h00000018; 
    validation_data[  179] = 'h00000088; 
    validation_data[  180] = 'h000003ce; 
    validation_data[  181] = 'h0000005a; 
    validation_data[  182] = 'h000003ef; 
    validation_data[  183] = 'h00000171; 
    validation_data[  184] = 'h00000134; 
    validation_data[  185] = 'h000002ac; 
    validation_data[  186] = 'h000003dc; 
    validation_data[  187] = 'h000000b1; 
    validation_data[  188] = 'h000002e6; 
    validation_data[  189] = 'h0000006e; 
    validation_data[  190] = 'h0000034d; 
    validation_data[  191] = 'h000001cb; 
    validation_data[  192] = 'h000000e2; 
    validation_data[  193] = 'h0000003e; 
    validation_data[  194] = 'h0000035d; 
    validation_data[  195] = 'h0000008e; 
    validation_data[  196] = 'h00000289; 
    validation_data[  197] = 'h000003bb; 
    validation_data[  198] = 'h000003a3; 
    validation_data[  199] = 'h00000391; 
    validation_data[  200] = 'h00000395; 
    validation_data[  201] = 'h000003be; 
    validation_data[  202] = 'h0000028d; 
    validation_data[  203] = 'h0000022c; 
    validation_data[  204] = 'h000003ca; 
    validation_data[  205] = 'h000002e2; 
    validation_data[  206] = 'h0000000e; 
    validation_data[  207] = 'h000002ac; 
    validation_data[  208] = 'h0000031f; 
    validation_data[  209] = 'h00000105; 
    validation_data[  210] = 'h000001c1; 
    validation_data[  211] = 'h00000361; 
    validation_data[  212] = 'h000002bd; 
    validation_data[  213] = 'h00000314; 
    validation_data[  214] = 'h0000026d; 
    validation_data[  215] = 'h0000025d; 
    validation_data[  216] = 'h000003ea; 
    validation_data[  217] = 'h0000005c; 
    validation_data[  218] = 'h000001f1; 
    validation_data[  219] = 'h000002fb; 
    validation_data[  220] = 'h000002d1; 
    validation_data[  221] = 'h000001c0; 
    validation_data[  222] = 'h00000344; 
    validation_data[  223] = 'h000002fa; 
    validation_data[  224] = 'h0000022e; 
    validation_data[  225] = 'h000000d3; 
    validation_data[  226] = 'h00000271; 
    validation_data[  227] = 'h00000383; 
    validation_data[  228] = 'h00000050; 
    validation_data[  229] = 'h000002d6; 
    validation_data[  230] = 'h0000014f; 
    validation_data[  231] = 'h000003be; 
    validation_data[  232] = 'h00000198; 
    validation_data[  233] = 'h000000fe; 
    validation_data[  234] = 'h0000036a; 
    validation_data[  235] = 'h00000088; 
    validation_data[  236] = 'h000001b2; 
    validation_data[  237] = 'h00000147; 
    validation_data[  238] = 'h000001a7; 
    validation_data[  239] = 'h000001ca; 
    validation_data[  240] = 'h00000045; 
    validation_data[  241] = 'h00000391; 
    validation_data[  242] = 'h0000030d; 
    validation_data[  243] = 'h000001b3; 
    validation_data[  244] = 'h0000018c; 
    validation_data[  245] = 'h0000033e; 
    validation_data[  246] = 'h00000114; 
    validation_data[  247] = 'h0000036e; 
    validation_data[  248] = 'h000001e3; 
    validation_data[  249] = 'h00000177; 
    validation_data[  250] = 'h000000a0; 
    validation_data[  251] = 'h00000153; 
    validation_data[  252] = 'h0000039f; 
    validation_data[  253] = 'h000000ce; 
    validation_data[  254] = 'h00000291; 
    validation_data[  255] = 'h000002c5; 

end


reg clk = 1'b1, rst = 1'b1;
initial #4 rst = 1'b0;
always  #1 clk = ~clk;

wire  miss;
wire [31:0] rd_data;
reg  [31:0] index = 0, wr_data = 0, addr = 0;
reg  rd_req = 1'b0, wr_req = 1'b0;
reg rd_req_ff = 1'b0, miss_ff = 1'b0;
reg [31:0] validation_count = 0;

always @ (posedge clk or posedge rst)
    if(rst) begin
        rd_req_ff <= 1'b0;
        miss_ff   <= 1'b0;
    end else begin
        rd_req_ff <= rd_req;
        miss_ff   <= miss;
    end

always @ (posedge clk or posedge rst)
    if(rst) begin
        validation_count <= 0;
    end else begin
        if(validation_count>=`DATA_COUNT) begin
            validation_count <= 'hffffffff;
        end else if(rd_req_ff && (index>(4*`DATA_COUNT))) begin
            if(~miss_ff) begin
                if(validation_data[validation_count]==rd_data)
                    validation_count <= validation_count+1;
                else
                    validation_count <= 0;
            end
        end else begin
            validation_count <= 0;
        end
    end

always @ (posedge clk or posedge rst)
    if(rst) begin
        index   <= 0;
        wr_data <= 0;
        addr    <= 0;
        rd_req  <= 1'b0;
        wr_req  <= 1'b0;
    end else begin
        if(~miss) begin
            if(index<`RDWR_COUNT) begin
                if(wr_cycle[index]) begin
                    rd_req  <= 1'b0;
                    wr_req  <= 1'b1;
                end else if(rd_cycle[index]) begin
                    wr_data <= 0;
                    rd_req  <= 1'b1;
                    wr_req  <= 1'b0;
                end else begin
                    wr_data <= 0;
                    rd_req  <= 1'b0;
                    wr_req  <= 1'b0;
                end
                wr_data <= wr_data_rom[index];
                addr    <= addr_rom[index];
                index <= index + 1;
            end else begin
                wr_data <= 0;
                addr    <= 0;
                rd_req  <= 1'b0;
                wr_req  <= 1'b0;
            end
        end
    end

cache #(
    .LINE_ADDR_LEN  ( 3             ),
    .SET_ADDR_LEN   ( 2             ),
    .TAG_ADDR_LEN   ( 12            ),
    .WAY_CNT        ( 3             )
) cache_test_instance (
    .clk            ( clk           ),
    .rst            ( rst           ),
    .miss           ( miss          ),
    .addr           ( addr          ),
    .rd_req         ( rd_req        ),
    .rd_data        ( rd_data       ),
    .wr_req         ( wr_req        ),
    .wr_data        ( wr_data       )
);

endmodule

